
//------> ./softmax_sysc_Connections_OutBlockingless_dma_info_tcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_sysc_Connections_OutBlockingless_dma_info_tcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_sysc_Connections_OutBlockingless_dma_info_tcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue Jun  9 12:18:22 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core
    (
  this_val, this_rdy, this_msg, m_index_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [66:0] this_msg;
  input [31:0] m_index_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire [31:0] m_index_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [24:0] m_index_slc_m_index_31_7_psp_lpi_1_dfm;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  reg reg_C_35_1_reg_32;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd32)) m_index_rsci (
      .dat(m_index_rsc_dat),
      .idat(m_index_rsci_idat)
    );
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 #(.rscid(32'sd45),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 #(.rscid(32'sd50)) ccs_ccore_done_synci
      (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign this_msg = {1'b0 , ({{1{reg_C_35_1_reg_32}}, reg_C_35_1_reg_32}) , 24'b000000000000000000000000
      , reg_C_35_1_reg_32 , 7'b0000000 , m_index_slc_m_index_31_7_psp_lpi_1_dfm ,
      7'b0000000};
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_val <= 1'b0;
    end
    else if ( or_4_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      reg_C_35_1_reg_32 <= 1'b0;
    end
    else if ( (~((~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1) | this_rdy)) | ccs_ccore_start_rsci_idat
        ) begin
      reg_C_35_1_reg_32 <= 1'b1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      m_index_slc_m_index_31_7_psp_lpi_1_dfm <= 25'b0000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      m_index_slc_m_index_31_7_psp_lpi_1_dfm <= m_index_rsci_idat[31:7];
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_index_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  input this_rdy;
  output [66:0] this_msg;
  input [31:0] m_index_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core_inst (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_index_rsc_dat(m_index_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_sysc_Connections_InBlockingless_dma_data_tcomma_Connections_SYN_PORTgreater_Pop_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./softmax_sysc_Connections_InBlockingless_dma_data_tcomma_Connections_SYN_PORTgreater_Pop_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_sysc_Connections_InBlockingless_dma_data_tcomma_Connections_SYN_PORTgreater_Pop_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_sysc_Connections_InBlockingless_dma_data_tcomma_Connections_SYN_PORTgreater_Pop.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue Jun  9 12:18:26 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_Connections_InBlocking_dma_data_t_Connections_SYN_PORT_Pop_core
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_Connections_InBlocking_dma_data_t_Connections_SYN_PORT_Pop_core
    (
  this_val, this_rdy, this_msg, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [63:0] this_msg;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_2_cse;
  wire this_rdy_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [63:0] nl_return_rsci_d;
  assign nl_return_rsci_d = this_msg;
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_val;
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_mgc_out_dreg_v2 #(.rscid(32'sd4),
  .width(32'sd64)) return_rsci (
      .d(nl_return_rsci_d[63:0]),
      .z(return_rsc_z)
    );
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 #(.rscid(32'sd44),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 #(.rscid(32'sd49)) ccs_ccore_done_synci
      (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign or_2_cse = ccs_ccore_start_rsci_idat | (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_val));
  assign this_rdy_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_val
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_rdy <= 1'b0;
    end
    else if ( or_2_cse | this_rdy_mx0c1 ) begin
      this_rdy <= ~ this_rdy_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_2_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_dma_data_t_Connections_SYN_PORT_Pop
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_Connections_InBlocking_dma_data_t_Connections_SYN_PORT_Pop (
  this_val, this_rdy, this_msg, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  input this_val;
  output this_rdy;
  input [63:0] this_msg;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_Connections_InBlocking_dma_data_t_Connections_SYN_PORT_Pop_core
      Connections_InBlocking_dma_data_t_Connections_SYN_PORT_Pop_core_inst (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_sysc_handshake_t_req_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_sysc_handshake_t_req_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_sysc_handshake_t_req.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue Jun  9 12:18:24 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_handshake_t_req_core
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_handshake_t_req_core (
  this_req_req, this_ack_ack, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld, ccs_MIO_clk,
      ccs_MIO_srst
);
  output this_req_req;
  reg this_req_req;
  input this_ack_ack;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg do_asn_mdf_sva_st_1;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_st_2;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = do_asn_mdf_sva_st_1 & io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_st_2;
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 #(.rscid(32'sd43),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 #(.rscid(32'sd48)) ccs_ccore_done_synci
      (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_req_req <= 1'b0;
      do_asn_mdf_sva_st_1 <= 1'b0;
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_st_2 <= 1'b0;
    end
    else begin
      this_req_req <= io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_ack_ack;
      do_asn_mdf_sva_st_1 <= this_ack_ack;
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= ccs_ccore_start_rsci_idat |
          (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_ack_ack));
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_st_2 <= io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    handshake_t_req
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_handshake_t_req (
  this_req_req, this_ack_ack, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld, ccs_MIO_clk,
      ccs_MIO_srst
);
  output this_req_req;
  input this_ack_ack;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_handshake_t_req_core handshake_t_req_core_inst (
      .this_req_req(this_req_req),
      .this_ack_ack(this_ack_ack),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_sysc_mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_sysc_mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./softmax_sysc_mgc_in_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_sysc_mgc_in_sync_v2 (vd, vz);
    parameter valid = 1;

    output vd;
    input  vz;

    wire   vd;

    assign vd = vz;

endmodule



//------> ./softmax_sysc_handshake_t_ack_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_sysc_handshake_t_ack_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_sysc_handshake_t_ack.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue Jun  9 12:18:23 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_handshake_t_ack_core
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_handshake_t_ack_core (
  this_req_req, this_ack_ack, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld, ccs_MIO_clk,
      ccs_MIO_srst
);
  input this_req_req;
  output this_ack_ack;
  reg this_ack_ack;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire asn_ccs_ccore_done_synci_ivld_and_cse;
  wire this_ack_ack_mx0c1;


  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 #(.rscid(32'sd42),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 #(.rscid(32'sd47)) ccs_ccore_done_synci
      (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(asn_ccs_ccore_done_synci_ivld_and_cse)
    );
  assign asn_ccs_ccore_done_synci_ivld_and_cse = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_req_req;
  assign this_ack_ack_mx0c1 = asn_ccs_ccore_done_synci_ivld_and_cse & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_ack_ack <= 1'b0;
    end
    else if ( (((~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1) | this_req_req) &
        ccs_ccore_start_rsci_idat) | this_ack_ack_mx0c1 ) begin
      this_ack_ack <= ~ this_ack_ack_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( ~(io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_req_req)) )
        begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    handshake_t_ack
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_handshake_t_ack (
  this_req_req, this_ack_ack, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld, ccs_MIO_clk,
      ccs_MIO_srst
);
  input this_req_req;
  output this_ack_ack;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_handshake_t_ack_core handshake_t_ack_core_inst (
      .this_req_req(this_req_req),
      .this_ack_ack(this_ack_ack),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_sysc_mgc_mul_pipe_beh.v 
//
// File:      $Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v
//
// BASELINE:  Catapult-C version 2006b.63
// MODIFIED:  2007-04-03, tnagler
//
// Note: this file uses Verilog2001 features;
//       please enable Verilog2001 in the flow!

module esp_acc_softmax_sysc_mgc_mul_pipe (a, b, clk, en, a_rst, s_rst, z);

    // Parameters:
    parameter integer width_a = 32'd4;  // input a bit width
    parameter         signd_a =  1'b1;  // input a type (1=signed, 0=unsigned)
    parameter integer width_b = 32'd4;  // input b bit width
    parameter         signd_b =  1'b1;  // input b type (1=signed, 0=unsigned)
    parameter integer width_z = 32'd8;  // result bit width (= width_a + width_b)
    parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
    parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
    parameter    a_rst_active =  1'b1;  // unused
    parameter    s_rst_active =  1'b1;  // unused
    parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
    parameter integer n_inreg = 32'd0;  // number of input registers

    localparam integer width_ab = width_a + width_b;  // multiplier result width
    localparam integer n_inreg_min = (n_inreg > 1) ? (n_inreg-1) : 0; // for Synopsys DC

    // I/O ports:
    input  [width_a-1:0] a;      // input A
    input  [width_b-1:0] b;      // input B
    input                clk;    // clock
    input                en;     // enable
    input                a_rst;  // async reset (unused)
    input                s_rst;  // sync reset (unused)
    output [width_z-1:0] z;      // output


    // Input registers:

    wire [width_a-1:0] a_f;
    wire [width_b-1:0] b_f;

    integer i;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(negedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i];
                    b_reg[i+1] <= b_reg[i];
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    else
    begin: POS_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(posedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i];
                    b_reg[i+1] <= b_reg[i];
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    endgenerate


    // Output:
    wire [width_z-1:0]  xz;

    function signed [width_z-1:0] conv_signed;
      input signed [width_ab-1:0] res;
      conv_signed = res[width_z-1:0];
    endfunction

    generate
      wire signed [width_ab-1:0] res;
      if ( (signd_a == 1'b1) && (signd_b == 1'b1) )
      begin: SIGNED_AB
              assign res = $signed(a_f) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b1) && (signd_b == 1'b0) )
      begin: SIGNED_A
              assign res = $signed(a_f) * $signed({1'b0, b_f});
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b0) && (signd_b == 1'b1) )
      begin: SIGNED_B
              assign res = $signed({1'b0,a_f}) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else
      begin: UNSIGNED_AB
              assign res = a_f * b_f;
	      assign xz = res[width_z-1:0];
      end
    endgenerate


    // Output registers:

    reg  [width_z-1:0] reg_array[stages-2:0];
    wire [width_z-1:0] z;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE2
        always @(negedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz;
                else
                    reg_array[i] <= reg_array[i-1];
    end
    else
    begin: POS_EDGE2
        always @(posedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz;
                else
                    reg_array[i] <= reg_array[i-1];
    end
    endgenerate

    assign z = reg_array[stages-2];
endmodule

//------> ./softmax_sysc_mgc_shift_br_beh_v5.v 
module esp_acc_softmax_sysc_mgc_shift_br_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_s(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_s(a,s,1'b0);
     end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshr_u

   //Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction

endmodule

//------> ./softmax_sysc_mgc_shift_bl_beh_v5.v 
module esp_acc_softmax_sysc_mgc_shift_bl_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate if ( signd_a )
   begin: SGNED
     assign z = fshl_s(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
     assign z = fshl_s(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

endmodule

//------> ./softmax_sysc_mgc_shift_l_beh_v5.v 
module esp_acc_softmax_sysc_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./softmax_sysc_leading_sign_74_0.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue Jun  9 12:18:25 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_74_0
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_leading_sign_74_0 (
  mantissa, rtn
);
  input [73:0] mantissa;
  output [6:0] rtn;


  // Interconnect Declarations
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_24;
  wire c_h_1_27;
  wire c_h_1_28;
  wire c_h_1_29;
  wire c_h_1_30;
  wire c_h_1_33;
  wire c_h_1_34;
  wire c_h_1_35;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc;

  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_1_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_292_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_2_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_or_2_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_nor_nl;

  // Interconnect Declarations for Component Instantiations
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2
      = ~((mantissa[71:70]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1
      = ~((mantissa[73:72]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1
      = ~((mantissa[69:68]!=2'b00));
  assign c_h_1_2 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3
      = (mantissa[67:66]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2
      = ~((mantissa[63:62]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1
      = ~((mantissa[65:64]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1
      = ~((mantissa[61:60]!=2'b00));
  assign c_h_1_5 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4
      = (mantissa[59:58]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1
      & c_h_1_5;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2
      = ~((mantissa[55:54]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1
      = ~((mantissa[57:56]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1
      = ~((mantissa[53:52]!=2'b00));
  assign c_h_1_9 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3
      = (mantissa[51:50]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2
      = ~((mantissa[47:46]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1
      = ~((mantissa[49:48]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1
      = ~((mantissa[45:44]!=2'b00));
  assign c_h_1_12 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5
      = (mantissa[43:42]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1
      & c_h_1_12 & c_h_1_13;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2
      = ~((mantissa[39:38]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1
      = ~((mantissa[41:40]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1
      = ~((mantissa[37:36]!=2'b00));
  assign c_h_1_17 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3
      = (mantissa[35:34]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2
      = ~((mantissa[31:30]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1
      = ~((mantissa[33:32]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1
      = ~((mantissa[29:28]!=2'b00));
  assign c_h_1_20 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4
      = (mantissa[27:26]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1
      & c_h_1_20;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2
      = ~((mantissa[23:22]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1
      = ~((mantissa[25:24]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1
      = ~((mantissa[21:20]!=2'b00));
  assign c_h_1_24 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3
      = (mantissa[19:18]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2
      = ~((mantissa[15:14]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1
      = ~((mantissa[17:16]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1
      = ~((mantissa[13:12]!=2'b00));
  assign c_h_1_27 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2;
  assign c_h_1_28 = c_h_1_24 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3;
  assign c_h_1_29 = c_h_1_21 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_30 = c_h_1_14 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6
      = (mantissa[11:10]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1
      & c_h_1_27 & c_h_1_28 & c_h_1_29;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2
      = ~((mantissa[7:6]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1
      = ~((mantissa[9:8]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1
      = ~((mantissa[5:4]!=2'b00));
  assign c_h_1_33 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3
      = (mantissa[3:2]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1;
  assign c_h_1_34 = c_h_1_33 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3;
  assign c_h_1_35 = c_h_1_30 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc
      = (mantissa[1:0]==2'b00) & c_h_1_34 & c_h_1_35;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_nl
      = c_h_1_30 & (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6);
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_1_nl
      = c_h_1_14 & (c_h_1_29 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5))
      & (~ c_h_1_35);
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_292_nl
      = c_h_1_6 & (c_h_1_13 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4))
      & (~((~(c_h_1_21 & (c_h_1_28 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4))))
      & c_h_1_30)) & (c_h_1_34 | (~ c_h_1_35));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_2_nl
      = c_h_1_2 & (c_h_1_5 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3))
      & (~((~(c_h_1_9 & (c_h_1_12 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~((~(c_h_1_17 & (c_h_1_20 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3))
      & (~((~(c_h_1_24 & (c_h_1_27 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3))))
      & c_h_1_29)))) & c_h_1_30)) & (~((~(c_h_1_33 & (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3)))
      & c_h_1_35));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_or_2_nl
      = (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2))))
      & c_h_1_21)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2))))
      & c_h_1_28)))) & c_h_1_29)))) & c_h_1_30)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2))
      & (~ c_h_1_34))) & c_h_1_35))) | ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_nor_nl
      = ~((mantissa[73]) | (~((mantissa[72:71]!=2'b01))) | (((mantissa[69]) | (~((mantissa[68:67]!=2'b01))))
      & c_h_1_2) | ((~((~((mantissa[65]) | (~((mantissa[64:63]!=2'b01))))) & (~(((mantissa[61])
      | (~((mantissa[60:59]!=2'b01)))) & c_h_1_5)))) & c_h_1_6) | ((~((~((mantissa[57])
      | (~((mantissa[56:55]!=2'b01))))) & (~(((mantissa[53]) | (~((mantissa[52:51]!=2'b01))))
      & c_h_1_9)) & (~((~((~((mantissa[49]) | (~((mantissa[48:47]!=2'b01))))) & (~(((mantissa[45])
      | (~((mantissa[44:43]!=2'b01)))) & c_h_1_12)))) & c_h_1_13)))) & c_h_1_14)
      | ((~((~((mantissa[41]) | (~((mantissa[40:39]!=2'b01))))) & (~(((mantissa[37])
      | (~((mantissa[36:35]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[33]) | (~((mantissa[32:31]!=2'b01)))))
      & (~(((mantissa[29]) | (~((mantissa[28:27]!=2'b01)))) & c_h_1_20)))) & c_h_1_21))
      & (~((~((~((mantissa[25]) | (~((mantissa[24:23]!=2'b01))))) & (~(((mantissa[21])
      | (~((mantissa[20:19]!=2'b01)))) & c_h_1_24)) & (~((~((~((mantissa[17]) | (~((mantissa[16:15]!=2'b01)))))
      & (~(((mantissa[13]) | (~((mantissa[12:11]!=2'b01)))) & c_h_1_27)))) & c_h_1_28))))
      & c_h_1_29)))) & c_h_1_30) | ((~((~((mantissa[9]) | (~((mantissa[8:7]!=2'b01)))))
      & (~(((mantissa[5]) | (~((mantissa[4:3]!=2'b01)))) & c_h_1_33)) & (~((mantissa[1])
      & c_h_1_34)))) & c_h_1_35) | ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc);
  assign rtn = {c_h_1_35 , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_1_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_292_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_2_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_or_2_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_nor_nl};
endmodule




//------> /opt/cad/catapult/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 
  
)( clk,clken,d,q,radr,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" *)
  reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block"
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./softmax_sysc_Connections_OutBlockingless_dma_data_tcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_sysc_Connections_OutBlockingless_dma_data_tcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_sysc_Connections_OutBlockingless_dma_data_tcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue Jun  9 12:18:21 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_Connections_OutBlocking_dma_data_t_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_Connections_OutBlocking_dma_data_t_Connections_SYN_PORT_Push_core
    (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [63:0] this_msg;
  input [63:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire [63:0] m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [31:0] m_slc_m_31_0_psp_lpi_1_dfm;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  reg reg_C_32_11011110101011011011111011101111_1_reg_30;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd64)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 #(.rscid(32'sd41),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 #(.rscid(32'sd46)) ccs_ccore_done_synci
      (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign this_msg = signext_64_63({reg_C_32_11011110101011011011111011101111_1_reg_30
      , 1'b0 , ({{3{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , reg_C_32_11011110101011011011111011101111_1_reg_30 , 1'b0 , reg_C_32_11011110101011011011111011101111_1_reg_30
      , 1'b0 , ({{1{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{1{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{4{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{2{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{3{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , m_slc_m_31_0_psp_lpi_1_dfm});
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_val <= 1'b0;
    end
    else if ( or_4_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      reg_C_32_11011110101011011011111011101111_1_reg_30 <= 1'b0;
    end
    else if ( (~((~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1) | this_rdy)) | ccs_ccore_start_rsci_idat
        ) begin
      reg_C_32_11011110101011011011111011101111_1_reg_30 <= 1'b1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      m_slc_m_31_0_psp_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      m_slc_m_31_0_psp_lpi_1_dfm <= m_rsci_idat[31:0];
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end

  function automatic [63:0] signext_64_63;
    input [62:0] vector;
  begin
    signext_64_63= {{1{vector[62]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_dma_data_t_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_Connections_OutBlocking_dma_data_t_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  input this_rdy;
  output [63:0] this_msg;
  input [63:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_Connections_OutBlocking_dma_data_t_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_dma_data_t_Connections_SYN_PORT_Push_core_inst (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_rsc_dat(m_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_sysc.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue Jun  9 12:18:55 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysczjlBRut_cns_bctl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysczjlBRut_cns_bctl (
  clk, rst, plm_out_cns_wadr_nsoftmax_sysc_compute_inst, plm_out_cns_d_nsoftmax_sysc_compute_inst,
      plm_out_cns_we_nsoftmax_sysc_compute_inst, plm_out_cns_req_vz_nsoftmax_sysc_compute_inst,
      plm_out_cns_we_nsoftmax_sysc_compute_inst_buz, plm_out_cns_radr_nsoftmax_sysc_store_inst,
      plm_out_cns_q_nsoftmax_sysc_store_inst, plm_out_cns_req_vz_nsoftmax_sysc_store_inst,
      plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud, plm_out_cns_rls_lz_nsoftmax_sysc_compute_inst_bud,
      plm_out_cns_rls_lz_nsoftmax_sysc_store_inst_bud, plm_out_cns_S0, plm_out_cns_R0,
      plm_out_cns_S1, plm_out_cns_R1, plm_out_cns_d_shi0, plm_out_cns_d_shi1, plm_out_cns_q_sho0,
      plm_out_cns_q_sho1, plm_out_cns_radr_shi0, plm_out_cns_radr_shi1, plm_out_cns_wadr_shi0,
      plm_out_cns_wadr_shi1, plm_out_cns_we_shi0, plm_out_cns_we_shi1, plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_pff,
      plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud_pff, plm_out_cns_S0_pff
);
  input clk;
  input rst;
  input [6:0] plm_out_cns_wadr_nsoftmax_sysc_compute_inst;
  input [31:0] plm_out_cns_d_nsoftmax_sysc_compute_inst;
  input plm_out_cns_we_nsoftmax_sysc_compute_inst;
  output plm_out_cns_req_vz_nsoftmax_sysc_compute_inst;
  input plm_out_cns_we_nsoftmax_sysc_compute_inst_buz;
  input [6:0] plm_out_cns_radr_nsoftmax_sysc_store_inst;
  output [31:0] plm_out_cns_q_nsoftmax_sysc_store_inst;
  output plm_out_cns_req_vz_nsoftmax_sysc_store_inst;
  output plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud;
  input plm_out_cns_rls_lz_nsoftmax_sysc_compute_inst_bud;
  input plm_out_cns_rls_lz_nsoftmax_sysc_store_inst_bud;
  output plm_out_cns_S0;
  input plm_out_cns_R0;
  output plm_out_cns_S1;
  input plm_out_cns_R1;
  output [31:0] plm_out_cns_d_shi0;
  output [31:0] plm_out_cns_d_shi1;
  input [31:0] plm_out_cns_q_sho0;
  input [31:0] plm_out_cns_q_sho1;
  output [6:0] plm_out_cns_radr_shi0;
  output [6:0] plm_out_cns_radr_shi1;
  output [6:0] plm_out_cns_wadr_shi0;
  output [6:0] plm_out_cns_wadr_shi1;
  output plm_out_cns_we_shi0;
  output plm_out_cns_we_shi1;
  input plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_pff;
  output plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud_pff;
  output plm_out_cns_S0_pff;


  // Interconnect Declarations
  reg plm_out_cns_we_nsoftmax_sysc_compute_inst_buy;
  wire plm_out_cns_PC0;
  reg plm_out_cns_ppidx;
  reg [1:0] plm_out_cns_ppown;
  wire plm_out_cns_PC1;
  reg plm_out_cns_ppidx_1;
  reg [1:0] plm_out_cns_ppown_1;
  wire [1:0] plm_out_acc_rmff;
  wire [3:0] nl_plm_out_acc_rmff;
  wire plm_out_xor_rmff;
  wire [1:0] plm_out_acc_1_rmff;
  wire [3:0] nl_plm_out_acc_1_rmff;


  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_req_vz_nsoftmax_sysc_compute_inst = plm_out_cns_R0;
  assign plm_out_cns_req_vz_nsoftmax_sysc_store_inst = plm_out_cns_R1;
  assign plm_out_xor_rmff = plm_out_cns_ppidx ^ plm_out_cns_PC0;
  assign nl_plm_out_acc_rmff = plm_out_cns_ppown + conv_u2u_1_2(plm_out_cns_PC0)
      + conv_s2u_1_2(plm_out_cns_PC1);
  assign plm_out_acc_rmff = nl_plm_out_acc_rmff[1:0];
  assign plm_out_cns_PC0 = plm_out_cns_S0 & plm_out_cns_rls_lz_nsoftmax_sysc_compute_inst_bud;
  assign nl_plm_out_acc_1_rmff = plm_out_cns_ppown_1 + conv_u2u_1_2(plm_out_cns_PC1)
      + conv_s2u_1_2(plm_out_cns_PC0);
  assign plm_out_acc_1_rmff = nl_plm_out_acc_1_rmff[1:0];
  assign plm_out_cns_PC1 = ((plm_out_cns_ppown_1!=2'b00)) & plm_out_cns_rls_lz_nsoftmax_sysc_store_inst_bud;
  assign plm_out_cns_q_nsoftmax_sysc_store_inst = MUX_v_32_2_2(plm_out_cns_q_sho0,
      plm_out_cns_q_sho1, plm_out_cns_ppidx_1);
  assign plm_out_cns_d_shi0 = plm_out_cns_d_nsoftmax_sysc_compute_inst;
  assign plm_out_cns_radr_shi0 = plm_out_cns_radr_nsoftmax_sysc_store_inst;
  assign plm_out_cns_wadr_shi0 = plm_out_cns_wadr_nsoftmax_sysc_compute_inst;
  assign plm_out_cns_we_shi0 = plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_pff
      & plm_out_cns_S0_pff & (~ plm_out_xor_rmff);
  assign plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud = plm_out_cns_we_nsoftmax_sysc_compute_inst_buy;
  assign plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud_pff = plm_out_cns_we_nsoftmax_sysc_compute_inst;
  assign plm_out_cns_S0 = ~((plm_out_cns_ppown==2'b10));
  assign plm_out_cns_S0_pff = ~((plm_out_acc_rmff==2'b10));
  assign plm_out_cns_d_shi1 = plm_out_cns_d_nsoftmax_sysc_compute_inst;
  assign plm_out_cns_radr_shi1 = plm_out_cns_radr_nsoftmax_sysc_store_inst;
  assign plm_out_cns_wadr_shi1 = plm_out_cns_wadr_nsoftmax_sysc_compute_inst;
  assign plm_out_cns_we_shi1 = plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_pff
      & plm_out_cns_S0_pff & plm_out_xor_rmff;
  assign plm_out_cns_S1 = (plm_out_acc_1_rmff!=2'b00);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cns_we_nsoftmax_sysc_compute_inst_buy <= 1'b0;
      plm_out_cns_ppidx <= 1'b0;
      plm_out_cns_ppown <= 2'b00;
      plm_out_cns_ppidx_1 <= 1'b0;
      plm_out_cns_ppown_1 <= 2'b00;
    end
    else begin
      plm_out_cns_we_nsoftmax_sysc_compute_inst_buy <= plm_out_cns_we_nsoftmax_sysc_compute_inst;
      plm_out_cns_ppidx <= plm_out_xor_rmff;
      plm_out_cns_ppown <= plm_out_acc_rmff;
      plm_out_cns_ppidx_1 <= plm_out_cns_ppidx_1 ^ plm_out_cns_PC1;
      plm_out_cns_ppown_1 <= plm_out_acc_1_rmff;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_plm_in_cns_bctl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_plm_in_cns_bctl (
  clk, rst, plm_in_cns_wadr_nsoftmax_sysc_load_inst, plm_in_cns_d_nsoftmax_sysc_load_inst,
      plm_in_cns_we_nsoftmax_sysc_load_inst, plm_in_cns_req_vz_nsoftmax_sysc_load_inst,
      plm_in_cns_radr_nsoftmax_sysc_compute_inst, plm_in_cns_q_nsoftmax_sysc_compute_inst,
      plm_in_cns_req_vz_nsoftmax_sysc_compute_inst, plm_out_cns_we_nsoftmax_sysc_compute_inst_buz,
      plm_in_cns_rls_lz_nsoftmax_sysc_load_inst_bud, plm_in_cns_rls_lz_nsoftmax_sysc_compute_inst_bud,
      plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud, plm_out_cns_rls_lz_nsoftmax_sysc_compute_inst_bud,
      plm_in_cns_S0, plm_in_cns_R0, plm_in_cns_S1, plm_in_cns_R1, plm_in_cns_d_shi0,
      plm_in_cns_d_shi1, plm_in_cns_q_sho0, plm_in_cns_q_sho1, plm_in_cns_radr_shi0,
      plm_in_cns_radr_shi1, plm_in_cns_wadr_shi0, plm_in_cns_wadr_shi1, plm_in_cns_we_shi0,
      plm_in_cns_we_shi1, plm_in_cns_S0_pff, plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_pff,
      plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud_pff
);
  input clk;
  input rst;
  input [6:0] plm_in_cns_wadr_nsoftmax_sysc_load_inst;
  input [31:0] plm_in_cns_d_nsoftmax_sysc_load_inst;
  input plm_in_cns_we_nsoftmax_sysc_load_inst;
  output plm_in_cns_req_vz_nsoftmax_sysc_load_inst;
  input [6:0] plm_in_cns_radr_nsoftmax_sysc_compute_inst;
  output [31:0] plm_in_cns_q_nsoftmax_sysc_compute_inst;
  output plm_in_cns_req_vz_nsoftmax_sysc_compute_inst;
  output plm_out_cns_we_nsoftmax_sysc_compute_inst_buz;
  input plm_in_cns_rls_lz_nsoftmax_sysc_load_inst_bud;
  input plm_in_cns_rls_lz_nsoftmax_sysc_compute_inst_bud;
  input plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud;
  input plm_out_cns_rls_lz_nsoftmax_sysc_compute_inst_bud;
  output plm_in_cns_S0;
  input plm_in_cns_R0;
  output plm_in_cns_S1;
  input plm_in_cns_R1;
  output [31:0] plm_in_cns_d_shi0;
  output [31:0] plm_in_cns_d_shi1;
  input [31:0] plm_in_cns_q_sho0;
  input [31:0] plm_in_cns_q_sho1;
  output [6:0] plm_in_cns_radr_shi0;
  output [6:0] plm_in_cns_radr_shi1;
  output [6:0] plm_in_cns_wadr_shi0;
  output [6:0] plm_in_cns_wadr_shi1;
  output plm_in_cns_we_shi0;
  output plm_in_cns_we_shi1;
  output plm_in_cns_S0_pff;
  output plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_pff;
  input plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud_pff;


  // Interconnect Declarations
  wire plm_in_cns_PC0;
  reg plm_in_cns_ppidx;
  reg [1:0] plm_in_cns_ppown;
  wire plm_in_cns_PC1;
  reg plm_in_cns_ppidx_1;
  reg [1:0] plm_in_cns_ppown_1;
  wire [1:0] plm_in_acc_rmff;
  wire [3:0] nl_plm_in_acc_rmff;
  wire plm_in_xor_rmff;
  wire [1:0] plm_in_acc_1_rmff;
  wire [3:0] nl_plm_in_acc_1_rmff;


  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_req_vz_nsoftmax_sysc_load_inst = plm_in_cns_R0;
  assign plm_in_cns_req_vz_nsoftmax_sysc_compute_inst = plm_in_cns_R1;
  assign plm_in_xor_rmff = plm_in_cns_ppidx ^ plm_in_cns_PC0;
  assign nl_plm_in_acc_rmff = plm_in_cns_ppown + conv_u2u_1_2(plm_in_cns_PC0) + conv_s2u_1_2(plm_in_cns_PC1);
  assign plm_in_acc_rmff = nl_plm_in_acc_rmff[1:0];
  assign plm_in_cns_PC0 = plm_in_cns_S0 & plm_in_cns_rls_lz_nsoftmax_sysc_load_inst_bud;
  assign nl_plm_in_acc_1_rmff = plm_in_cns_ppown_1 + conv_u2u_1_2(plm_in_cns_PC1)
      + conv_s2u_1_2(plm_in_cns_PC0);
  assign plm_in_acc_1_rmff = nl_plm_in_acc_1_rmff[1:0];
  assign plm_in_cns_PC1 = ((plm_in_cns_ppown_1!=2'b00)) & plm_in_cns_rls_lz_nsoftmax_sysc_compute_inst_bud;
  assign plm_in_cns_q_nsoftmax_sysc_compute_inst = MUX_v_32_2_2(plm_in_cns_q_sho0,
      plm_in_cns_q_sho1, plm_in_cns_ppidx_1);
  assign plm_in_cns_d_shi0 = plm_in_cns_d_nsoftmax_sysc_load_inst;
  assign plm_in_cns_radr_shi0 = plm_in_cns_radr_nsoftmax_sysc_compute_inst;
  assign plm_in_cns_wadr_shi0 = plm_in_cns_wadr_nsoftmax_sysc_load_inst;
  assign plm_in_cns_we_shi0 = plm_in_cns_we_nsoftmax_sysc_load_inst & plm_in_cns_S0_pff
      & (~ plm_in_xor_rmff);
  assign plm_in_cns_S0 = ~((plm_in_cns_ppown==2'b10));
  assign plm_in_cns_S0_pff = ~((plm_in_acc_rmff==2'b10));
  assign plm_in_cns_d_shi1 = plm_in_cns_d_nsoftmax_sysc_load_inst;
  assign plm_in_cns_radr_shi1 = plm_in_cns_radr_nsoftmax_sysc_compute_inst;
  assign plm_in_cns_wadr_shi1 = plm_in_cns_wadr_nsoftmax_sysc_load_inst;
  assign plm_in_cns_we_shi1 = plm_in_cns_we_nsoftmax_sysc_load_inst & plm_in_cns_S0_pff
      & plm_in_xor_rmff;
  assign plm_out_cns_we_nsoftmax_sysc_compute_inst_buz = plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud;
  assign plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_pff = plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud_pff;
  assign plm_in_cns_S1 = (plm_in_acc_1_rmff!=2'b00);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cns_ppidx <= 1'b0;
      plm_in_cns_ppown <= 2'b00;
      plm_in_cns_ppidx_1 <= 1'b0;
      plm_in_cns_ppown_1 <= 2'b00;
    end
    else begin
      plm_in_cns_ppidx <= plm_in_xor_rmff;
      plm_in_cns_ppown <= plm_in_acc_rmff;
      plm_in_cns_ppidx_1 <= plm_in_cns_ppidx_1 ^ plm_in_cns_PC1;
      plm_in_cns_ppown_1 <= plm_in_acc_1_rmff;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_unreg_hier
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_unreg_hier (
  in_0, out_0
);
  input in_0;
  output out_0;



  // Interconnect Declarations for Component Instantiations 
  assign out_0 = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_7_32_128_128_32_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_7_32_128_128_32_1_gen
    (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [6:0] radr;
  output [31:0] q_d;
  input [6:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_store_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_store_fsm (
  clk, rst, store_wen, fsm_output, WAIT_FOR_CONFIG_LOOP_C_0_tr0, STORE_BATCH_LOOP_C_0_tr0
);
  input clk;
  input rst;
  input store_wen;
  output [6:0] fsm_output;
  reg [6:0] fsm_output;
  input WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  input STORE_BATCH_LOOP_C_0_tr0;


  // FSM State Type Declaration for esp_acc_softmax_sysc_softmax_sysc_store_store_store_fsm_1
  parameter
    WAIT_FOR_CONFIG_LOOP_C_0 = 3'd0,
    STORE_BATCH_LOOP_C_0 = 3'd1,
    store_rlp_C_0 = 3'd2,
    store_rlp_C_1 = 3'd3,
    store_rlp_C_2 = 3'd4,
    store_rlp_C_3 = 3'd5,
    PROCESS_DONE_LOOP_C_0 = 3'd6;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_softmax_sysc_softmax_sysc_store_store_store_fsm_1
    case (state_var)
      STORE_BATCH_LOOP_C_0 : begin
        fsm_output = 7'b0000010;
        if ( STORE_BATCH_LOOP_C_0_tr0 ) begin
          state_var_NS = STORE_BATCH_LOOP_C_0;
        end
        else begin
          state_var_NS = store_rlp_C_0;
        end
      end
      store_rlp_C_0 : begin
        fsm_output = 7'b0000100;
        state_var_NS = store_rlp_C_1;
      end
      store_rlp_C_1 : begin
        fsm_output = 7'b0001000;
        state_var_NS = store_rlp_C_2;
      end
      store_rlp_C_2 : begin
        fsm_output = 7'b0010000;
        state_var_NS = store_rlp_C_3;
      end
      store_rlp_C_3 : begin
        fsm_output = 7'b0100000;
        state_var_NS = PROCESS_DONE_LOOP_C_0;
      end
      PROCESS_DONE_LOOP_C_0 : begin
        fsm_output = 7'b1000000;
        state_var_NS = PROCESS_DONE_LOOP_C_0;
      end
      // WAIT_FOR_CONFIG_LOOP_C_0
      default : begin
        fsm_output = 7'b0000001;
        if ( WAIT_FOR_CONFIG_LOOP_C_0_tr0 ) begin
          state_var_NS = WAIT_FOR_CONFIG_LOOP_C_0;
        end
        else begin
          state_var_NS = STORE_BATCH_LOOP_C_0;
        end
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= WAIT_FOR_CONFIG_LOOP_C_0;
    end
    else if ( store_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_staller
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_staller (
  clk, rst, store_wen, store_wten, output_ready_ack_mioi_wen_comp, dma_write_ctrl_Push_mioi_wen_comp,
      dma_write_chnl_Push_mioi_wen_comp, plm_out_cns_req_obj_wen_comp
);
  input clk;
  input rst;
  output store_wen;
  output store_wten;
  input output_ready_ack_mioi_wen_comp;
  input dma_write_ctrl_Push_mioi_wen_comp;
  input dma_write_chnl_Push_mioi_wen_comp;
  input plm_out_cns_req_obj_wen_comp;


  // Interconnect Declarations
  reg store_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign store_wen = output_ready_ack_mioi_wen_comp & dma_write_ctrl_Push_mioi_wen_comp
      & dma_write_chnl_Push_mioi_wen_comp & plm_out_cns_req_obj_wen_comp;
  assign store_wten = store_wten_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      store_wten_reg <= 1'b0;
    end
    else begin
      store_wten_reg <= ~ store_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_req_obj_plm_out_cns_req_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_req_obj_plm_out_cns_req_wait_dp
    (
  clk, rst, plm_out_cns_req_obj_oswt_unreg, plm_out_cns_req_obj_bawt, plm_out_cns_req_obj_wen_comp,
      plm_out_cns_req_obj_biwt, plm_out_cns_req_obj_bdwt, plm_out_cns_req_obj_bcwt
);
  input clk;
  input rst;
  input plm_out_cns_req_obj_oswt_unreg;
  output plm_out_cns_req_obj_bawt;
  output plm_out_cns_req_obj_wen_comp;
  input plm_out_cns_req_obj_biwt;
  input plm_out_cns_req_obj_bdwt;
  output plm_out_cns_req_obj_bcwt;
  reg plm_out_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_req_obj_bawt = plm_out_cns_req_obj_biwt | plm_out_cns_req_obj_bcwt;
  assign plm_out_cns_req_obj_wen_comp = (~ plm_out_cns_req_obj_oswt_unreg) | plm_out_cns_req_obj_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cns_req_obj_bcwt <= 1'b0;
    end
    else begin
      plm_out_cns_req_obj_bcwt <= ~((~(plm_out_cns_req_obj_bcwt | plm_out_cns_req_obj_biwt))
          | plm_out_cns_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl
    (
  store_wen, plm_out_cns_req_obj_oswt_unreg, plm_out_cns_req_obj_iswt0, plm_out_cns_req_obj_vd,
      plm_out_cns_req_obj_biwt, plm_out_cns_req_obj_bdwt, plm_out_cns_req_obj_bcwt
);
  input store_wen;
  input plm_out_cns_req_obj_oswt_unreg;
  input plm_out_cns_req_obj_iswt0;
  input plm_out_cns_req_obj_vd;
  output plm_out_cns_req_obj_biwt;
  output plm_out_cns_req_obj_bdwt;
  input plm_out_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_req_obj_bdwt = plm_out_cns_req_obj_oswt_unreg & store_wen;
  assign plm_out_cns_req_obj_biwt = plm_out_cns_req_obj_iswt0 & (~ plm_out_cns_req_obj_bcwt)
      & plm_out_cns_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_rls_obj_plm_out_cns_rls_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_rls_obj_plm_out_cns_rls_wait_dp
    (
  clk, rst, plm_out_cns_rls_obj_bawt, plm_out_cns_rls_obj_biwt, plm_out_cns_rls_obj_bdwt
);
  input clk;
  input rst;
  output plm_out_cns_rls_obj_bawt;
  input plm_out_cns_rls_obj_biwt;
  input plm_out_cns_rls_obj_bdwt;


  // Interconnect Declarations
  reg plm_out_cns_rls_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_rls_obj_bawt = plm_out_cns_rls_obj_biwt | plm_out_cns_rls_obj_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cns_rls_obj_bcwt <= 1'b0;
    end
    else begin
      plm_out_cns_rls_obj_bcwt <= ~((~(plm_out_cns_rls_obj_bcwt | plm_out_cns_rls_obj_biwt))
          | plm_out_cns_rls_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl
    (
  store_wen, store_wten, plm_out_cns_rls_obj_oswt_unreg, plm_out_cns_rls_obj_iswt0,
      plm_out_cns_rls_obj_biwt, plm_out_cns_rls_obj_bdwt
);
  input store_wen;
  input store_wten;
  input plm_out_cns_rls_obj_oswt_unreg;
  input plm_out_cns_rls_obj_iswt0;
  output plm_out_cns_rls_obj_biwt;
  output plm_out_cns_rls_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_rls_obj_bdwt = plm_out_cns_rls_obj_oswt_unreg & store_wen;
  assign plm_out_cns_rls_obj_biwt = (~ store_wten) & plm_out_cns_rls_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cnsi_1_plm_out_cns_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cnsi_1_plm_out_cns_wait_dp
    (
  clk, rst, plm_out_cnsi_q_d, plm_out_cnsi_bawt, plm_out_cnsi_q_d_mxwt, plm_out_cnsi_biwt,
      plm_out_cnsi_bdwt
);
  input clk;
  input rst;
  input [31:0] plm_out_cnsi_q_d;
  output plm_out_cnsi_bawt;
  output [31:0] plm_out_cnsi_q_d_mxwt;
  input plm_out_cnsi_biwt;
  input plm_out_cnsi_bdwt;


  // Interconnect Declarations
  reg plm_out_cnsi_bcwt;
  reg [31:0] plm_out_cnsi_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cnsi_bawt = plm_out_cnsi_biwt | plm_out_cnsi_bcwt;
  assign plm_out_cnsi_q_d_mxwt = MUX_v_32_2_2(plm_out_cnsi_q_d, plm_out_cnsi_q_d_bfwt,
      plm_out_cnsi_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cnsi_bcwt <= 1'b0;
    end
    else begin
      plm_out_cnsi_bcwt <= ~((~(plm_out_cnsi_bcwt | plm_out_cnsi_biwt)) | plm_out_cnsi_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( plm_out_cnsi_biwt ) begin
      plm_out_cnsi_q_d_bfwt <= plm_out_cnsi_q_d;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cnsi_1_plm_out_cns_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cnsi_1_plm_out_cns_wait_ctrl
    (
  store_wen, store_wten, plm_out_cnsi_oswt_unreg, plm_out_cnsi_iswt0, plm_out_cnsi_biwt,
      plm_out_cnsi_bdwt, plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_store_sct,
      plm_out_cnsi_iswt0_pff
);
  input store_wen;
  input store_wten;
  input plm_out_cnsi_oswt_unreg;
  input plm_out_cnsi_iswt0;
  output plm_out_cnsi_biwt;
  output plm_out_cnsi_bdwt;
  output plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_store_sct;
  input plm_out_cnsi_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cnsi_bdwt = plm_out_cnsi_oswt_unreg & store_wen;
  assign plm_out_cnsi_biwt = (~ store_wten) & plm_out_cnsi_iswt0;
  assign plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_store_sct = plm_out_cnsi_iswt0_pff
      & store_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp
    (
  clk, rst, dma_write_chnl_Push_mioi_oswt_unreg, dma_write_chnl_Push_mioi_bawt, dma_write_chnl_Push_mioi_wen_comp,
      dma_write_chnl_Push_mioi_biwt, dma_write_chnl_Push_mioi_bdwt
);
  input clk;
  input rst;
  input dma_write_chnl_Push_mioi_oswt_unreg;
  output dma_write_chnl_Push_mioi_bawt;
  output dma_write_chnl_Push_mioi_wen_comp;
  input dma_write_chnl_Push_mioi_biwt;
  input dma_write_chnl_Push_mioi_bdwt;


  // Interconnect Declarations
  reg dma_write_chnl_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_write_chnl_Push_mioi_bawt = dma_write_chnl_Push_mioi_biwt | dma_write_chnl_Push_mioi_bcwt;
  assign dma_write_chnl_Push_mioi_wen_comp = (~ dma_write_chnl_Push_mioi_oswt_unreg)
      | dma_write_chnl_Push_mioi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_chnl_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_write_chnl_Push_mioi_bcwt <= ~((~(dma_write_chnl_Push_mioi_bcwt | dma_write_chnl_Push_mioi_biwt))
          | dma_write_chnl_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl
    (
  clk, rst, store_wen, store_wten, dma_write_chnl_Push_mioi_oswt_unreg, dma_write_chnl_Push_mioi_iswt0,
      dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct, dma_write_chnl_Push_mioi_biwt,
      dma_write_chnl_Push_mioi_bdwt, dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_sct,
      dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld, dma_write_chnl_Push_mioi_iswt0_pff
);
  input clk;
  input rst;
  input store_wen;
  input store_wten;
  input dma_write_chnl_Push_mioi_oswt_unreg;
  input dma_write_chnl_Push_mioi_iswt0;
  input dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct;
  output dma_write_chnl_Push_mioi_biwt;
  output dma_write_chnl_Push_mioi_bdwt;
  output dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_sct;
  input dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld;
  input dma_write_chnl_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire dma_write_chnl_Push_mioi_ogwt;
  reg dma_write_chnl_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_write_chnl_Push_mioi_bdwt = dma_write_chnl_Push_mioi_oswt_unreg & store_wen;
  assign dma_write_chnl_Push_mioi_biwt = dma_write_chnl_Push_mioi_ogwt & dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld;
  assign dma_write_chnl_Push_mioi_ogwt = ((~ store_wten) & dma_write_chnl_Push_mioi_iswt0)
      | dma_write_chnl_Push_mioi_icwt;
  assign dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_sct = dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct
      & store_wen & dma_write_chnl_Push_mioi_iswt0_pff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_chnl_Push_mioi_icwt <= 1'b0;
    end
    else begin
      dma_write_chnl_Push_mioi_icwt <= dma_write_chnl_Push_mioi_ogwt & (~ dma_write_chnl_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp
    (
  clk, rst, dma_write_ctrl_Push_mioi_oswt_unreg, dma_write_ctrl_Push_mioi_bawt, dma_write_ctrl_Push_mioi_wen_comp,
      dma_write_ctrl_Push_mioi_biwt, dma_write_ctrl_Push_mioi_bdwt
);
  input clk;
  input rst;
  input dma_write_ctrl_Push_mioi_oswt_unreg;
  output dma_write_ctrl_Push_mioi_bawt;
  output dma_write_ctrl_Push_mioi_wen_comp;
  input dma_write_ctrl_Push_mioi_biwt;
  input dma_write_ctrl_Push_mioi_bdwt;


  // Interconnect Declarations
  reg dma_write_ctrl_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_write_ctrl_Push_mioi_bawt = dma_write_ctrl_Push_mioi_biwt | dma_write_ctrl_Push_mioi_bcwt;
  assign dma_write_ctrl_Push_mioi_wen_comp = (~ dma_write_ctrl_Push_mioi_oswt_unreg)
      | dma_write_ctrl_Push_mioi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_ctrl_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_write_ctrl_Push_mioi_bcwt <= ~((~(dma_write_ctrl_Push_mioi_bcwt | dma_write_ctrl_Push_mioi_biwt))
          | dma_write_ctrl_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl
    (
  clk, rst, store_wen, store_wten, dma_write_ctrl_Push_mioi_oswt_unreg, dma_write_ctrl_Push_mioi_iswt0,
      dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct, dma_write_ctrl_Push_mioi_biwt,
      dma_write_ctrl_Push_mioi_bdwt, dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_sct,
      dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld, dma_write_ctrl_Push_mioi_iswt0_pff
);
  input clk;
  input rst;
  input store_wen;
  input store_wten;
  input dma_write_ctrl_Push_mioi_oswt_unreg;
  input dma_write_ctrl_Push_mioi_iswt0;
  input dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct;
  output dma_write_ctrl_Push_mioi_biwt;
  output dma_write_ctrl_Push_mioi_bdwt;
  output dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_sct;
  input dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  input dma_write_ctrl_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire dma_write_ctrl_Push_mioi_ogwt;
  reg dma_write_ctrl_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_write_ctrl_Push_mioi_bdwt = dma_write_ctrl_Push_mioi_oswt_unreg & store_wen;
  assign dma_write_ctrl_Push_mioi_biwt = dma_write_ctrl_Push_mioi_ogwt & dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  assign dma_write_ctrl_Push_mioi_ogwt = ((~ store_wten) & dma_write_ctrl_Push_mioi_iswt0)
      | dma_write_ctrl_Push_mioi_icwt;
  assign dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_sct = dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct
      & store_wen & dma_write_ctrl_Push_mioi_iswt0_pff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_ctrl_Push_mioi_icwt <= 1'b0;
    end
    else begin
      dma_write_ctrl_Push_mioi_icwt <= dma_write_ctrl_Push_mioi_ogwt & (~ dma_write_ctrl_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_output_ready_ack_mioi_output_ready_ack_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_output_ready_ack_mioi_output_ready_ack_mio_wait_dp
    (
  clk, rst, output_ready_ack_mioi_oswt_unreg, output_ready_ack_mioi_bawt, output_ready_ack_mioi_wen_comp,
      output_ready_ack_mioi_biwt, output_ready_ack_mioi_bdwt
);
  input clk;
  input rst;
  input output_ready_ack_mioi_oswt_unreg;
  output output_ready_ack_mioi_bawt;
  output output_ready_ack_mioi_wen_comp;
  input output_ready_ack_mioi_biwt;
  input output_ready_ack_mioi_bdwt;


  // Interconnect Declarations
  reg output_ready_ack_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign output_ready_ack_mioi_bawt = output_ready_ack_mioi_biwt | output_ready_ack_mioi_bcwt;
  assign output_ready_ack_mioi_wen_comp = (~ output_ready_ack_mioi_oswt_unreg) |
      output_ready_ack_mioi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      output_ready_ack_mioi_bcwt <= 1'b0;
    end
    else begin
      output_ready_ack_mioi_bcwt <= ~((~(output_ready_ack_mioi_bcwt | output_ready_ack_mioi_biwt))
          | output_ready_ack_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_output_ready_ack_mioi_output_ready_ack_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_output_ready_ack_mioi_output_ready_ack_mio_wait_ctrl
    (
  clk, rst, store_wen, output_ready_ack_mioi_oswt_unreg, output_ready_ack_mioi_iswt0,
      store_wten, output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_psct, output_ready_ack_mioi_biwt,
      output_ready_ack_mioi_bdwt, output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_sct,
      output_ready_ack_mioi_ccs_ccore_done_sync_vld, output_ready_ack_mioi_iswt0_pff
);
  input clk;
  input rst;
  input store_wen;
  input output_ready_ack_mioi_oswt_unreg;
  input output_ready_ack_mioi_iswt0;
  input store_wten;
  input output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_psct;
  output output_ready_ack_mioi_biwt;
  output output_ready_ack_mioi_bdwt;
  output output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_sct;
  input output_ready_ack_mioi_ccs_ccore_done_sync_vld;
  input output_ready_ack_mioi_iswt0_pff;


  // Interconnect Declarations
  wire output_ready_ack_mioi_ogwt;
  reg output_ready_ack_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign output_ready_ack_mioi_bdwt = output_ready_ack_mioi_oswt_unreg & store_wen;
  assign output_ready_ack_mioi_biwt = output_ready_ack_mioi_ogwt & output_ready_ack_mioi_ccs_ccore_done_sync_vld;
  assign output_ready_ack_mioi_ogwt = ((~ store_wten) & output_ready_ack_mioi_iswt0)
      | output_ready_ack_mioi_icwt;
  assign output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_sct = output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_psct
      & store_wen & output_ready_ack_mioi_iswt0_pff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      output_ready_ack_mioi_icwt <= 1'b0;
    end
    else begin
      output_ready_ack_mioi_icwt <= output_ready_ack_mioi_ogwt & (~ output_ready_ack_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_35_7_32_128_128_32_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_35_7_32_128_128_32_1_gen
    (
  we, d, wadr, d_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [31:0] d;
  output [6:0] wadr;
  input [31:0] d_d;
  input [6:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_7_32_128_128_32_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_7_32_128_128_32_1_gen
    (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [6:0] radr;
  output [31:0] q_d;
  input [6:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_17_7_67_128_128_67_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_17_7_67_128_128_67_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [66:0] q;
  output [6:0] radr;
  output we;
  output [66:0] d;
  output [6:0] wadr;
  input clken_d;
  input [66:0] d_d;
  output [66:0] q_d;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_compute_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_compute_fsm (
  clk, rst, compute_wen, fsm_output, WAIT_FOR_CONFIG_LOOP_C_0_tr0, COMPUTE_BATCH_LOOP_C_0_tr0
);
  input clk;
  input rst;
  input compute_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;
  input WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  input COMPUTE_BATCH_LOOP_C_0_tr0;


  // FSM State Type Declaration for esp_acc_softmax_sysc_softmax_sysc_compute_compute_compute_fsm_1
  parameter
    WAIT_FOR_CONFIG_LOOP_C_0 = 2'd0,
    COMPUTE_BATCH_LOOP_C_0 = 2'd1,
    PROCESS_DONE_LOOP_C_0 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_softmax_sysc_softmax_sysc_compute_compute_compute_fsm_1
    case (state_var)
      COMPUTE_BATCH_LOOP_C_0 : begin
        fsm_output = 3'b010;
        if ( COMPUTE_BATCH_LOOP_C_0_tr0 ) begin
          state_var_NS = COMPUTE_BATCH_LOOP_C_0;
        end
        else begin
          state_var_NS = PROCESS_DONE_LOOP_C_0;
        end
      end
      PROCESS_DONE_LOOP_C_0 : begin
        fsm_output = 3'b100;
        state_var_NS = PROCESS_DONE_LOOP_C_0;
      end
      // WAIT_FOR_CONFIG_LOOP_C_0
      default : begin
        fsm_output = 3'b001;
        if ( WAIT_FOR_CONFIG_LOOP_C_0_tr0 ) begin
          state_var_NS = WAIT_FOR_CONFIG_LOOP_C_0;
        end
        else begin
          state_var_NS = COMPUTE_BATCH_LOOP_C_0;
        end
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= WAIT_FOR_CONFIG_LOOP_C_0;
    end
    else if ( compute_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_staller
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_staller (
  clk, rst, compute_wen, compute_wten, input_ready_ack_mioi_wen_comp, output_ready_req_mioi_wen_comp,
      plm_in_cns_req_obj_wen_comp, plm_out_cns_req_obj_wen_comp
);
  input clk;
  input rst;
  output compute_wen;
  output compute_wten;
  input input_ready_ack_mioi_wen_comp;
  input output_ready_req_mioi_wen_comp;
  input plm_in_cns_req_obj_wen_comp;
  input plm_out_cns_req_obj_wen_comp;


  // Interconnect Declarations
  reg compute_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign compute_wen = input_ready_ack_mioi_wen_comp & output_ready_req_mioi_wen_comp
      & plm_in_cns_req_obj_wen_comp & plm_out_cns_req_obj_wen_comp;
  assign compute_wten = compute_wten_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      compute_wten_reg <= 1'b0;
    end
    else begin
      compute_wten_reg <= ~ compute_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_req_obj_plm_out_cns_req_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_req_obj_plm_out_cns_req_wait_dp
    (
  clk, rst, plm_out_cns_req_obj_oswt_unreg, plm_out_cns_req_obj_bawt, plm_out_cns_req_obj_wen_comp,
      plm_out_cns_req_obj_biwt, plm_out_cns_req_obj_bdwt, plm_out_cns_req_obj_bcwt
);
  input clk;
  input rst;
  input plm_out_cns_req_obj_oswt_unreg;
  output plm_out_cns_req_obj_bawt;
  output plm_out_cns_req_obj_wen_comp;
  input plm_out_cns_req_obj_biwt;
  input plm_out_cns_req_obj_bdwt;
  output plm_out_cns_req_obj_bcwt;
  reg plm_out_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_req_obj_bawt = plm_out_cns_req_obj_biwt | plm_out_cns_req_obj_bcwt;
  assign plm_out_cns_req_obj_wen_comp = (~ plm_out_cns_req_obj_oswt_unreg) | plm_out_cns_req_obj_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cns_req_obj_bcwt <= 1'b0;
    end
    else begin
      plm_out_cns_req_obj_bcwt <= ~((~(plm_out_cns_req_obj_bcwt | plm_out_cns_req_obj_biwt))
          | plm_out_cns_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl
    (
  compute_wen, plm_out_cns_req_obj_oswt_unreg, plm_out_cns_req_obj_iswt0, plm_out_cns_req_obj_vd,
      plm_out_cns_req_obj_biwt, plm_out_cns_req_obj_bdwt, plm_out_cns_req_obj_bcwt
);
  input compute_wen;
  input plm_out_cns_req_obj_oswt_unreg;
  input plm_out_cns_req_obj_iswt0;
  input plm_out_cns_req_obj_vd;
  output plm_out_cns_req_obj_biwt;
  output plm_out_cns_req_obj_bdwt;
  input plm_out_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_req_obj_bdwt = plm_out_cns_req_obj_oswt_unreg & compute_wen;
  assign plm_out_cns_req_obj_biwt = plm_out_cns_req_obj_iswt0 & (~ plm_out_cns_req_obj_bcwt)
      & plm_out_cns_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_req_obj_plm_in_cns_req_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_req_obj_plm_in_cns_req_wait_dp
    (
  clk, rst, plm_in_cns_req_obj_oswt_unreg, plm_in_cns_req_obj_bawt, plm_in_cns_req_obj_wen_comp,
      plm_in_cns_req_obj_biwt, plm_in_cns_req_obj_bdwt, plm_in_cns_req_obj_bcwt
);
  input clk;
  input rst;
  input plm_in_cns_req_obj_oswt_unreg;
  output plm_in_cns_req_obj_bawt;
  output plm_in_cns_req_obj_wen_comp;
  input plm_in_cns_req_obj_biwt;
  input plm_in_cns_req_obj_bdwt;
  output plm_in_cns_req_obj_bcwt;
  reg plm_in_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_req_obj_bawt = plm_in_cns_req_obj_biwt | plm_in_cns_req_obj_bcwt;
  assign plm_in_cns_req_obj_wen_comp = (~ plm_in_cns_req_obj_oswt_unreg) | plm_in_cns_req_obj_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cns_req_obj_bcwt <= 1'b0;
    end
    else begin
      plm_in_cns_req_obj_bcwt <= ~((~(plm_in_cns_req_obj_bcwt | plm_in_cns_req_obj_biwt))
          | plm_in_cns_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl
    (
  compute_wen, plm_in_cns_req_obj_oswt_unreg, plm_in_cns_req_obj_iswt0, plm_in_cns_req_obj_vd,
      plm_in_cns_req_obj_biwt, plm_in_cns_req_obj_bdwt, plm_in_cns_req_obj_bcwt
);
  input compute_wen;
  input plm_in_cns_req_obj_oswt_unreg;
  input plm_in_cns_req_obj_iswt0;
  input plm_in_cns_req_obj_vd;
  output plm_in_cns_req_obj_biwt;
  output plm_in_cns_req_obj_bdwt;
  input plm_in_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_req_obj_bdwt = plm_in_cns_req_obj_oswt_unreg & compute_wen;
  assign plm_in_cns_req_obj_biwt = plm_in_cns_req_obj_iswt0 & (~ plm_in_cns_req_obj_bcwt)
      & plm_in_cns_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_rls_obj_plm_in_cns_rls_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_rls_obj_plm_in_cns_rls_wait_dp
    (
  clk, rst, plm_in_cns_rls_obj_bawt, plm_in_cns_rls_obj_biwt, plm_in_cns_rls_obj_bdwt
);
  input clk;
  input rst;
  output plm_in_cns_rls_obj_bawt;
  input plm_in_cns_rls_obj_biwt;
  input plm_in_cns_rls_obj_bdwt;


  // Interconnect Declarations
  reg plm_in_cns_rls_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_rls_obj_bawt = plm_in_cns_rls_obj_biwt | plm_in_cns_rls_obj_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cns_rls_obj_bcwt <= 1'b0;
    end
    else begin
      plm_in_cns_rls_obj_bcwt <= ~((~(plm_in_cns_rls_obj_bcwt | plm_in_cns_rls_obj_biwt))
          | plm_in_cns_rls_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl
    (
  compute_wen, compute_wten, plm_in_cns_rls_obj_oswt_unreg, plm_in_cns_rls_obj_iswt0,
      plm_in_cns_rls_obj_biwt, plm_in_cns_rls_obj_bdwt
);
  input compute_wen;
  input compute_wten;
  input plm_in_cns_rls_obj_oswt_unreg;
  input plm_in_cns_rls_obj_iswt0;
  output plm_in_cns_rls_obj_biwt;
  output plm_in_cns_rls_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_rls_obj_bdwt = plm_in_cns_rls_obj_oswt_unreg & compute_wen;
  assign plm_in_cns_rls_obj_biwt = (~ compute_wten) & plm_in_cns_rls_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_dp
    (
  clk, rst, CALC_SOFTMAX_LOOP_mul_cmp_bawt, CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt, CALC_SOFTMAX_LOOP_mul_cmp_biwt,
      CALC_SOFTMAX_LOOP_mul_cmp_bdwt, CALC_SOFTMAX_LOOP_mul_cmp_z
);
  input clk;
  input rst;
  output CALC_SOFTMAX_LOOP_mul_cmp_bawt;
  output [31:0] CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt;
  input CALC_SOFTMAX_LOOP_mul_cmp_biwt;
  input CALC_SOFTMAX_LOOP_mul_cmp_bdwt;
  input [94:0] CALC_SOFTMAX_LOOP_mul_cmp_z;


  // Interconnect Declarations
  reg [1:0] CALC_SOFTMAX_LOOP_mul_cmp_bcwt;
  wire [2:0] nl_CALC_SOFTMAX_LOOP_mul_cmp_bcwt;
  reg [31:0] CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_2_94_63;
  reg [31:0] CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_1_94_63;
  reg [31:0] CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_94_63;

  wire[1:0] CALC_SOFTMAX_LOOP_acc_1_nl;
  wire[2:0] nl_CALC_SOFTMAX_LOOP_acc_1_nl;
  wire[1:0] CALC_SOFTMAX_LOOP_acc_2_nl;
  wire[2:0] nl_CALC_SOFTMAX_LOOP_acc_2_nl;

  // Interconnect Declarations for Component Instantiations 
  assign CALC_SOFTMAX_LOOP_mul_cmp_bawt = CALC_SOFTMAX_LOOP_mul_cmp_biwt | (CALC_SOFTMAX_LOOP_mul_cmp_bcwt!=2'b00);
  assign CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt = MUX_v_32_4_2((CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]),
      CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_94_63, CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_1_94_63,
      CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_2_94_63, CALC_SOFTMAX_LOOP_mul_cmp_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_mul_cmp_bcwt <= 2'b00;
    end
    else begin
      CALC_SOFTMAX_LOOP_mul_cmp_bcwt <= nl_CALC_SOFTMAX_LOOP_mul_cmp_bcwt[1:0];
    end
  end
  always @(posedge clk) begin
    if ( CALC_SOFTMAX_LOOP_mul_cmp_biwt ) begin
      CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_94_63 <= CALC_SOFTMAX_LOOP_mul_cmp_z[94:63];
      CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_1_94_63 <= CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_94_63;
      CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_2_94_63 <= CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_1_94_63;
    end
  end
  assign nl_CALC_SOFTMAX_LOOP_acc_1_nl = conv_u2u_1_2(CALC_SOFTMAX_LOOP_mul_cmp_biwt)
      + conv_u2u_1_2(~ CALC_SOFTMAX_LOOP_mul_cmp_bdwt);
  assign CALC_SOFTMAX_LOOP_acc_1_nl = nl_CALC_SOFTMAX_LOOP_acc_1_nl[1:0];
  assign nl_CALC_SOFTMAX_LOOP_acc_2_nl = CALC_SOFTMAX_LOOP_mul_cmp_bcwt + 2'b11;
  assign CALC_SOFTMAX_LOOP_acc_2_nl = nl_CALC_SOFTMAX_LOOP_acc_2_nl[1:0];
  assign nl_CALC_SOFTMAX_LOOP_mul_cmp_bcwt  = CALC_SOFTMAX_LOOP_acc_1_nl + CALC_SOFTMAX_LOOP_acc_2_nl;

  function automatic [31:0] MUX_v_32_4_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [31:0] input_3;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_32_4_2 = result;
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_ctrl
    (
  clk, rst, compute_wen, compute_wten, CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg, CALC_SOFTMAX_LOOP_mul_cmp_iswt2,
      CALC_SOFTMAX_LOOP_mul_cmp_biwt, CALC_SOFTMAX_LOOP_mul_cmp_bdwt
);
  input clk;
  input rst;
  input compute_wen;
  input compute_wten;
  input CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg;
  input CALC_SOFTMAX_LOOP_mul_cmp_iswt2;
  output CALC_SOFTMAX_LOOP_mul_cmp_biwt;
  output CALC_SOFTMAX_LOOP_mul_cmp_bdwt;


  // Interconnect Declarations
  reg CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt1;
  reg CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt0;
  reg [1:0] CALC_SOFTMAX_LOOP_mul_cmp_icwt;
  wire [2:0] nl_CALC_SOFTMAX_LOOP_mul_cmp_icwt;

  wire[1:0] CALC_SOFTMAX_LOOP_acc_2_nl;
  wire[2:0] nl_CALC_SOFTMAX_LOOP_acc_2_nl;
  wire[1:0] CALC_SOFTMAX_LOOP_acc_3_nl;
  wire[2:0] nl_CALC_SOFTMAX_LOOP_acc_3_nl;

  // Interconnect Declarations for Component Instantiations 
  assign CALC_SOFTMAX_LOOP_mul_cmp_bdwt = CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg &
      compute_wen;
  assign CALC_SOFTMAX_LOOP_mul_cmp_biwt = CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt0
      | (CALC_SOFTMAX_LOOP_mul_cmp_icwt!=2'b00);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt1 <= 1'b0;
      CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt0 <= 1'b0;
      CALC_SOFTMAX_LOOP_mul_cmp_icwt <= 2'b00;
    end
    else begin
      CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt1 <= (~ compute_wten)
          & CALC_SOFTMAX_LOOP_mul_cmp_iswt2;
      CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt0 <= CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt1;
      CALC_SOFTMAX_LOOP_mul_cmp_icwt <= nl_CALC_SOFTMAX_LOOP_mul_cmp_icwt[1:0];
    end
  end
  assign nl_CALC_SOFTMAX_LOOP_acc_2_nl = conv_u2u_1_2(CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt0)
      + conv_u2u_1_2(~ CALC_SOFTMAX_LOOP_mul_cmp_biwt);
  assign CALC_SOFTMAX_LOOP_acc_2_nl = nl_CALC_SOFTMAX_LOOP_acc_2_nl[1:0];
  assign nl_CALC_SOFTMAX_LOOP_acc_3_nl = CALC_SOFTMAX_LOOP_mul_cmp_icwt + 2'b11;
  assign CALC_SOFTMAX_LOOP_acc_3_nl = nl_CALC_SOFTMAX_LOOP_acc_3_nl[1:0];
  assign nl_CALC_SOFTMAX_LOOP_mul_cmp_icwt  = CALC_SOFTMAX_LOOP_acc_2_nl + CALC_SOFTMAX_LOOP_acc_3_nl;

  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_rls_obj_plm_out_cns_rls_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_rls_obj_plm_out_cns_rls_wait_dp
    (
  clk, rst, plm_out_cns_rls_obj_bawt, plm_out_cns_rls_obj_biwt, plm_out_cns_rls_obj_bdwt
);
  input clk;
  input rst;
  output plm_out_cns_rls_obj_bawt;
  input plm_out_cns_rls_obj_biwt;
  input plm_out_cns_rls_obj_bdwt;


  // Interconnect Declarations
  reg plm_out_cns_rls_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_rls_obj_bawt = plm_out_cns_rls_obj_biwt | plm_out_cns_rls_obj_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cns_rls_obj_bcwt <= 1'b0;
    end
    else begin
      plm_out_cns_rls_obj_bcwt <= ~((~(plm_out_cns_rls_obj_bcwt | plm_out_cns_rls_obj_biwt))
          | plm_out_cns_rls_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl
    (
  compute_wen, compute_wten, plm_out_cns_rls_obj_oswt_unreg, plm_out_cns_rls_obj_iswt0,
      plm_out_cns_rls_obj_biwt, plm_out_cns_rls_obj_bdwt
);
  input compute_wen;
  input compute_wten;
  input plm_out_cns_rls_obj_oswt_unreg;
  input plm_out_cns_rls_obj_iswt0;
  output plm_out_cns_rls_obj_biwt;
  output plm_out_cns_rls_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_rls_obj_bdwt = plm_out_cns_rls_obj_oswt_unreg & compute_wen;
  assign plm_out_cns_rls_obj_biwt = (~ compute_wten) & plm_out_cns_rls_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cnsi_1_plm_out_cns_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cnsi_1_plm_out_cns_wait_dp
    (
  clk, rst, plm_out_cnsi_bawt, plm_out_cnsi_biwt, plm_out_cnsi_bdwt
);
  input clk;
  input rst;
  output plm_out_cnsi_bawt;
  input plm_out_cnsi_biwt;
  input plm_out_cnsi_bdwt;


  // Interconnect Declarations
  reg plm_out_cnsi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cnsi_bawt = plm_out_cnsi_biwt | plm_out_cnsi_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cnsi_bcwt <= 1'b0;
    end
    else begin
      plm_out_cnsi_bcwt <= ~((~(plm_out_cnsi_bcwt | plm_out_cnsi_biwt)) | plm_out_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cnsi_1_plm_out_cns_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cnsi_1_plm_out_cns_wait_ctrl
    (
  compute_wen, compute_wten, plm_out_cnsi_oswt_unreg, plm_out_cnsi_iswt0, plm_out_cnsi_biwt,
      plm_out_cnsi_bdwt, plm_out_cnsi_we_d_compute_sct_pff, plm_out_cnsi_iswt0_pff
);
  input compute_wen;
  input compute_wten;
  input plm_out_cnsi_oswt_unreg;
  input plm_out_cnsi_iswt0;
  output plm_out_cnsi_biwt;
  output plm_out_cnsi_bdwt;
  output plm_out_cnsi_we_d_compute_sct_pff;
  input plm_out_cnsi_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cnsi_bdwt = plm_out_cnsi_oswt_unreg & compute_wen;
  assign plm_out_cnsi_biwt = (~ compute_wten) & plm_out_cnsi_iswt0;
  assign plm_out_cnsi_we_d_compute_sct_pff = plm_out_cnsi_iswt0_pff & compute_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cnsi_1_plm_in_cns_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cnsi_1_plm_in_cns_wait_dp
    (
  clk, rst, plm_in_cnsi_q_d, plm_in_cnsi_bawt, plm_in_cnsi_q_d_mxwt, plm_in_cnsi_biwt,
      plm_in_cnsi_bdwt
);
  input clk;
  input rst;
  input [31:0] plm_in_cnsi_q_d;
  output plm_in_cnsi_bawt;
  output [31:0] plm_in_cnsi_q_d_mxwt;
  input plm_in_cnsi_biwt;
  input plm_in_cnsi_bdwt;


  // Interconnect Declarations
  reg plm_in_cnsi_bcwt;
  reg [31:0] plm_in_cnsi_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cnsi_bawt = plm_in_cnsi_biwt | plm_in_cnsi_bcwt;
  assign plm_in_cnsi_q_d_mxwt = MUX_v_32_2_2(plm_in_cnsi_q_d, plm_in_cnsi_q_d_bfwt,
      plm_in_cnsi_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cnsi_bcwt <= 1'b0;
    end
    else begin
      plm_in_cnsi_bcwt <= ~((~(plm_in_cnsi_bcwt | plm_in_cnsi_biwt)) | plm_in_cnsi_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( plm_in_cnsi_biwt ) begin
      plm_in_cnsi_q_d_bfwt <= plm_in_cnsi_q_d;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cnsi_1_plm_in_cns_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cnsi_1_plm_in_cns_wait_ctrl
    (
  compute_wen, compute_wten, plm_in_cnsi_oswt_unreg, plm_in_cnsi_iswt0, plm_in_cnsi_biwt,
      plm_in_cnsi_bdwt, plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_compute_sct,
      plm_in_cnsi_iswt0_pff
);
  input compute_wen;
  input compute_wten;
  input plm_in_cnsi_oswt_unreg;
  input plm_in_cnsi_iswt0;
  output plm_in_cnsi_biwt;
  output plm_in_cnsi_bdwt;
  output plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_compute_sct;
  input plm_in_cnsi_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cnsi_bdwt = plm_in_cnsi_oswt_unreg & compute_wen;
  assign plm_in_cnsi_biwt = (~ compute_wten) & plm_in_cnsi_iswt0;
  assign plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_compute_sct = plm_in_cnsi_iswt0_pff
      & compute_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_output_ready_req_mioi_output_ready_req_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_output_ready_req_mioi_output_ready_req_mio_wait_dp
    (
  clk, rst, output_ready_req_mioi_oswt_unreg, output_ready_req_mioi_bawt, output_ready_req_mioi_wen_comp,
      output_ready_req_mioi_biwt, output_ready_req_mioi_bdwt
);
  input clk;
  input rst;
  input output_ready_req_mioi_oswt_unreg;
  output output_ready_req_mioi_bawt;
  output output_ready_req_mioi_wen_comp;
  input output_ready_req_mioi_biwt;
  input output_ready_req_mioi_bdwt;


  // Interconnect Declarations
  reg output_ready_req_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign output_ready_req_mioi_bawt = output_ready_req_mioi_biwt | output_ready_req_mioi_bcwt;
  assign output_ready_req_mioi_wen_comp = (~ output_ready_req_mioi_oswt_unreg) |
      output_ready_req_mioi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      output_ready_req_mioi_bcwt <= 1'b0;
    end
    else begin
      output_ready_req_mioi_bcwt <= ~((~(output_ready_req_mioi_bcwt | output_ready_req_mioi_biwt))
          | output_ready_req_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_output_ready_req_mioi_output_ready_req_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_output_ready_req_mioi_output_ready_req_mio_wait_ctrl
    (
  clk, rst, compute_wen, compute_wten, output_ready_req_mioi_oswt_unreg, output_ready_req_mioi_iswt0,
      output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_psct, output_ready_req_mioi_biwt,
      output_ready_req_mioi_bdwt, output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_sct,
      output_ready_req_mioi_ccs_ccore_done_sync_vld, output_ready_req_mioi_iswt0_pff
);
  input clk;
  input rst;
  input compute_wen;
  input compute_wten;
  input output_ready_req_mioi_oswt_unreg;
  input output_ready_req_mioi_iswt0;
  input output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_psct;
  output output_ready_req_mioi_biwt;
  output output_ready_req_mioi_bdwt;
  output output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_sct;
  input output_ready_req_mioi_ccs_ccore_done_sync_vld;
  input output_ready_req_mioi_iswt0_pff;


  // Interconnect Declarations
  wire output_ready_req_mioi_ogwt;
  reg output_ready_req_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign output_ready_req_mioi_bdwt = output_ready_req_mioi_oswt_unreg & compute_wen;
  assign output_ready_req_mioi_biwt = output_ready_req_mioi_ogwt & output_ready_req_mioi_ccs_ccore_done_sync_vld;
  assign output_ready_req_mioi_ogwt = ((~ compute_wten) & output_ready_req_mioi_iswt0)
      | output_ready_req_mioi_icwt;
  assign output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_sct = output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_psct
      & compute_wen & output_ready_req_mioi_iswt0_pff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      output_ready_req_mioi_icwt <= 1'b0;
    end
    else begin
      output_ready_req_mioi_icwt <= output_ready_req_mioi_ogwt & (~ output_ready_req_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_input_ready_ack_mioi_input_ready_ack_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_input_ready_ack_mioi_input_ready_ack_mio_wait_dp
    (
  clk, rst, input_ready_ack_mioi_oswt_unreg, input_ready_ack_mioi_bawt, input_ready_ack_mioi_wen_comp,
      input_ready_ack_mioi_biwt, input_ready_ack_mioi_bdwt
);
  input clk;
  input rst;
  input input_ready_ack_mioi_oswt_unreg;
  output input_ready_ack_mioi_bawt;
  output input_ready_ack_mioi_wen_comp;
  input input_ready_ack_mioi_biwt;
  input input_ready_ack_mioi_bdwt;


  // Interconnect Declarations
  reg input_ready_ack_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_ready_ack_mioi_bawt = input_ready_ack_mioi_biwt | input_ready_ack_mioi_bcwt;
  assign input_ready_ack_mioi_wen_comp = (~ input_ready_ack_mioi_oswt_unreg) | input_ready_ack_mioi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      input_ready_ack_mioi_bcwt <= 1'b0;
    end
    else begin
      input_ready_ack_mioi_bcwt <= ~((~(input_ready_ack_mioi_bcwt | input_ready_ack_mioi_biwt))
          | input_ready_ack_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_input_ready_ack_mioi_input_ready_ack_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_input_ready_ack_mioi_input_ready_ack_mio_wait_ctrl
    (
  clk, rst, compute_wen, compute_wten, input_ready_ack_mioi_oswt_unreg, input_ready_ack_mioi_iswt0,
      input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_psct, input_ready_ack_mioi_biwt,
      input_ready_ack_mioi_bdwt, input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_sct,
      input_ready_ack_mioi_ccs_ccore_done_sync_vld, input_ready_ack_mioi_iswt0_pff
);
  input clk;
  input rst;
  input compute_wen;
  input compute_wten;
  input input_ready_ack_mioi_oswt_unreg;
  input input_ready_ack_mioi_iswt0;
  input input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_psct;
  output input_ready_ack_mioi_biwt;
  output input_ready_ack_mioi_bdwt;
  output input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_sct;
  input input_ready_ack_mioi_ccs_ccore_done_sync_vld;
  input input_ready_ack_mioi_iswt0_pff;


  // Interconnect Declarations
  wire input_ready_ack_mioi_ogwt;
  reg input_ready_ack_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_ready_ack_mioi_bdwt = input_ready_ack_mioi_oswt_unreg & compute_wen;
  assign input_ready_ack_mioi_biwt = input_ready_ack_mioi_ogwt & input_ready_ack_mioi_ccs_ccore_done_sync_vld;
  assign input_ready_ack_mioi_ogwt = ((~ compute_wten) & input_ready_ack_mioi_iswt0)
      | input_ready_ack_mioi_icwt;
  assign input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_sct = input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_psct
      & compute_wen & input_ready_ack_mioi_iswt0_pff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      input_ready_ack_mioi_icwt <= 1'b0;
    end
    else begin
      input_ready_ack_mioi_icwt <= input_ready_ack_mioi_ogwt & (~ input_ready_ack_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_dp
    (
  clk, rst, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2
);
  input clk;
  input rst;
  input [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt;
  output [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2;


  // Interconnect Declarations
  reg ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt;
  reg ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt_1;
  reg [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt
      | ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt
      = MUX_v_67_2_2(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_bfwt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt_1);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt
          <= 1'b0;
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt_1
          <= 1'b0;
    end
    else begin
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt
          <= ~((~(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt
          | ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt))
          | ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt);
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt_1
          <= ~((~(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt_1
          | ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1))
          | ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2);
    end
  end
  always @(posedge clk) begin
    if ( ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1
        ) begin
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_bfwt
          <= ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d;
    end
  end

  function automatic [66:0] MUX_v_67_2_2;
    input [66:0] input_0;
    input [66:0] input_1;
    input [0:0] sel;
    reg [66:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_67_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_ctrl
    (
  compute_wen, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0,
      compute_wten, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_compute_sct,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_compute_sct_pff,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff
);
  input compute_wen;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0;
  input compute_wten;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_compute_sct;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_compute_sct_pff;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg
      & compute_wen;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt
      = (~ compute_wten) & ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1
      & compute_wen;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1
      = (~ compute_wten) & ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_compute_sct_pff
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff
      & compute_wen;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_compute_sct
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff
      & compute_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_33_7_32_128_128_32_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_33_7_32_128_128_32_1_gen
    (
  we, d, wadr, d_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [31:0] d;
  output [6:0] wadr;
  input [31:0] d_d;
  input [6:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_load_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_load_fsm (
  clk, rst, load_wen, fsm_output, WAIT_FOR_CONFIG_LOOP_C_0_tr0, LOAD_BATCH_LOOP_C_0_tr0
);
  input clk;
  input rst;
  input load_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;
  input WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  input LOAD_BATCH_LOOP_C_0_tr0;


  // FSM State Type Declaration for esp_acc_softmax_sysc_softmax_sysc_load_load_load_fsm_1
  parameter
    WAIT_FOR_CONFIG_LOOP_C_0 = 2'd0,
    LOAD_BATCH_LOOP_C_0 = 2'd1,
    PROCESS_DONE_LOOP_C_0 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_softmax_sysc_softmax_sysc_load_load_load_fsm_1
    case (state_var)
      LOAD_BATCH_LOOP_C_0 : begin
        fsm_output = 3'b010;
        if ( LOAD_BATCH_LOOP_C_0_tr0 ) begin
          state_var_NS = LOAD_BATCH_LOOP_C_0;
        end
        else begin
          state_var_NS = PROCESS_DONE_LOOP_C_0;
        end
      end
      PROCESS_DONE_LOOP_C_0 : begin
        fsm_output = 3'b100;
        state_var_NS = PROCESS_DONE_LOOP_C_0;
      end
      // WAIT_FOR_CONFIG_LOOP_C_0
      default : begin
        fsm_output = 3'b001;
        if ( WAIT_FOR_CONFIG_LOOP_C_0_tr0 ) begin
          state_var_NS = WAIT_FOR_CONFIG_LOOP_C_0;
        end
        else begin
          state_var_NS = LOAD_BATCH_LOOP_C_0;
        end
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= WAIT_FOR_CONFIG_LOOP_C_0;
    end
    else if ( load_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_staller
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_staller (
  clk, rst, load_wen, load_wten, dma_read_ctrl_Push_mioi_wen_comp, dma_read_chnl_Pop_mioi_wen_comp,
      input_ready_req_mioi_wen_comp, plm_in_cns_req_obj_wen_comp
);
  input clk;
  input rst;
  output load_wen;
  output load_wten;
  input dma_read_ctrl_Push_mioi_wen_comp;
  input dma_read_chnl_Pop_mioi_wen_comp;
  input input_ready_req_mioi_wen_comp;
  input plm_in_cns_req_obj_wen_comp;


  // Interconnect Declarations
  reg load_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign load_wen = dma_read_ctrl_Push_mioi_wen_comp & dma_read_chnl_Pop_mioi_wen_comp
      & input_ready_req_mioi_wen_comp & plm_in_cns_req_obj_wen_comp;
  assign load_wten = load_wten_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      load_wten_reg <= 1'b0;
    end
    else begin
      load_wten_reg <= ~ load_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_req_obj_plm_in_cns_req_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_req_obj_plm_in_cns_req_wait_dp
    (
  clk, rst, plm_in_cns_req_obj_oswt_unreg, plm_in_cns_req_obj_bawt, plm_in_cns_req_obj_wen_comp,
      plm_in_cns_req_obj_biwt, plm_in_cns_req_obj_bdwt, plm_in_cns_req_obj_bcwt
);
  input clk;
  input rst;
  input plm_in_cns_req_obj_oswt_unreg;
  output plm_in_cns_req_obj_bawt;
  output plm_in_cns_req_obj_wen_comp;
  input plm_in_cns_req_obj_biwt;
  input plm_in_cns_req_obj_bdwt;
  output plm_in_cns_req_obj_bcwt;
  reg plm_in_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_req_obj_bawt = plm_in_cns_req_obj_biwt | plm_in_cns_req_obj_bcwt;
  assign plm_in_cns_req_obj_wen_comp = (~ plm_in_cns_req_obj_oswt_unreg) | plm_in_cns_req_obj_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cns_req_obj_bcwt <= 1'b0;
    end
    else begin
      plm_in_cns_req_obj_bcwt <= ~((~(plm_in_cns_req_obj_bcwt | plm_in_cns_req_obj_biwt))
          | plm_in_cns_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl
    (
  load_wen, plm_in_cns_req_obj_oswt_unreg, plm_in_cns_req_obj_iswt0, plm_in_cns_req_obj_vd,
      plm_in_cns_req_obj_biwt, plm_in_cns_req_obj_bdwt, plm_in_cns_req_obj_bcwt
);
  input load_wen;
  input plm_in_cns_req_obj_oswt_unreg;
  input plm_in_cns_req_obj_iswt0;
  input plm_in_cns_req_obj_vd;
  output plm_in_cns_req_obj_biwt;
  output plm_in_cns_req_obj_bdwt;
  input plm_in_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_req_obj_bdwt = plm_in_cns_req_obj_oswt_unreg & load_wen;
  assign plm_in_cns_req_obj_biwt = plm_in_cns_req_obj_iswt0 & (~ plm_in_cns_req_obj_bcwt)
      & plm_in_cns_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_rls_obj_plm_in_cns_rls_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_rls_obj_plm_in_cns_rls_wait_dp
    (
  clk, rst, plm_in_cns_rls_obj_bawt, plm_in_cns_rls_obj_biwt, plm_in_cns_rls_obj_bdwt
);
  input clk;
  input rst;
  output plm_in_cns_rls_obj_bawt;
  input plm_in_cns_rls_obj_biwt;
  input plm_in_cns_rls_obj_bdwt;


  // Interconnect Declarations
  reg plm_in_cns_rls_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_rls_obj_bawt = plm_in_cns_rls_obj_biwt | plm_in_cns_rls_obj_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cns_rls_obj_bcwt <= 1'b0;
    end
    else begin
      plm_in_cns_rls_obj_bcwt <= ~((~(plm_in_cns_rls_obj_bcwt | plm_in_cns_rls_obj_biwt))
          | plm_in_cns_rls_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl
    (
  load_wen, load_wten, plm_in_cns_rls_obj_oswt_unreg, plm_in_cns_rls_obj_iswt0, plm_in_cns_rls_obj_biwt,
      plm_in_cns_rls_obj_bdwt
);
  input load_wen;
  input load_wten;
  input plm_in_cns_rls_obj_oswt_unreg;
  input plm_in_cns_rls_obj_iswt0;
  output plm_in_cns_rls_obj_biwt;
  output plm_in_cns_rls_obj_bdwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_rls_obj_bdwt = plm_in_cns_rls_obj_oswt_unreg & load_wen;
  assign plm_in_cns_rls_obj_biwt = (~ load_wten) & plm_in_cns_rls_obj_iswt0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cnsi_1_plm_in_cns_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cnsi_1_plm_in_cns_wait_dp
    (
  clk, rst, plm_in_cnsi_bawt, plm_in_cnsi_biwt, plm_in_cnsi_bdwt
);
  input clk;
  input rst;
  output plm_in_cnsi_bawt;
  input plm_in_cnsi_biwt;
  input plm_in_cnsi_bdwt;


  // Interconnect Declarations
  reg plm_in_cnsi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cnsi_bawt = plm_in_cnsi_biwt | plm_in_cnsi_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cnsi_bcwt <= 1'b0;
    end
    else begin
      plm_in_cnsi_bcwt <= ~((~(plm_in_cnsi_bcwt | plm_in_cnsi_biwt)) | plm_in_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cnsi_1_plm_in_cns_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cnsi_1_plm_in_cns_wait_ctrl
    (
  load_wen, load_wten, plm_in_cnsi_oswt_unreg, plm_in_cnsi_iswt0, plm_in_cnsi_biwt,
      plm_in_cnsi_bdwt, plm_in_cnsi_we_d_load_sct_pff, plm_in_cnsi_iswt0_pff
);
  input load_wen;
  input load_wten;
  input plm_in_cnsi_oswt_unreg;
  input plm_in_cnsi_iswt0;
  output plm_in_cnsi_biwt;
  output plm_in_cnsi_bdwt;
  output plm_in_cnsi_we_d_load_sct_pff;
  input plm_in_cnsi_iswt0_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cnsi_bdwt = plm_in_cnsi_oswt_unreg & load_wen;
  assign plm_in_cnsi_biwt = (~ load_wten) & plm_in_cnsi_iswt0;
  assign plm_in_cnsi_we_d_load_sct_pff = plm_in_cnsi_iswt0_pff & load_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_input_ready_req_mioi_input_ready_req_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_input_ready_req_mioi_input_ready_req_mio_wait_dp
    (
  clk, rst, input_ready_req_mioi_oswt_unreg, input_ready_req_mioi_bawt, input_ready_req_mioi_wen_comp,
      input_ready_req_mioi_biwt, input_ready_req_mioi_bdwt
);
  input clk;
  input rst;
  input input_ready_req_mioi_oswt_unreg;
  output input_ready_req_mioi_bawt;
  output input_ready_req_mioi_wen_comp;
  input input_ready_req_mioi_biwt;
  input input_ready_req_mioi_bdwt;


  // Interconnect Declarations
  reg input_ready_req_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_ready_req_mioi_bawt = input_ready_req_mioi_biwt | input_ready_req_mioi_bcwt;
  assign input_ready_req_mioi_wen_comp = (~ input_ready_req_mioi_oswt_unreg) | input_ready_req_mioi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      input_ready_req_mioi_bcwt <= 1'b0;
    end
    else begin
      input_ready_req_mioi_bcwt <= ~((~(input_ready_req_mioi_bcwt | input_ready_req_mioi_biwt))
          | input_ready_req_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_input_ready_req_mioi_input_ready_req_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_input_ready_req_mioi_input_ready_req_mio_wait_ctrl
    (
  clk, rst, load_wen, load_wten, input_ready_req_mioi_oswt_unreg, input_ready_req_mioi_iswt0,
      input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_psct, input_ready_req_mioi_biwt,
      input_ready_req_mioi_bdwt, input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_sct,
      input_ready_req_mioi_ccs_ccore_done_sync_vld, input_ready_req_mioi_iswt0_pff
);
  input clk;
  input rst;
  input load_wen;
  input load_wten;
  input input_ready_req_mioi_oswt_unreg;
  input input_ready_req_mioi_iswt0;
  input input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_psct;
  output input_ready_req_mioi_biwt;
  output input_ready_req_mioi_bdwt;
  output input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_sct;
  input input_ready_req_mioi_ccs_ccore_done_sync_vld;
  input input_ready_req_mioi_iswt0_pff;


  // Interconnect Declarations
  wire input_ready_req_mioi_ogwt;
  reg input_ready_req_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_ready_req_mioi_bdwt = input_ready_req_mioi_oswt_unreg & load_wen;
  assign input_ready_req_mioi_biwt = input_ready_req_mioi_ogwt & input_ready_req_mioi_ccs_ccore_done_sync_vld;
  assign input_ready_req_mioi_ogwt = ((~ load_wten) & input_ready_req_mioi_iswt0)
      | input_ready_req_mioi_icwt;
  assign input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_sct = input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_psct
      & load_wen & input_ready_req_mioi_iswt0_pff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      input_ready_req_mioi_icwt <= 1'b0;
    end
    else begin
      input_ready_req_mioi_icwt <= input_ready_req_mioi_ogwt & (~ input_ready_req_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp
    (
  clk, rst, dma_read_chnl_Pop_mioi_oswt_unreg, dma_read_chnl_Pop_mioi_bawt, dma_read_chnl_Pop_mioi_wen_comp,
      dma_read_chnl_Pop_mioi_return_rsc_z_mxwt, dma_read_chnl_Pop_mioi_return_rsc_z,
      dma_read_chnl_Pop_mioi_biwt, dma_read_chnl_Pop_mioi_bdwt
);
  input clk;
  input rst;
  input dma_read_chnl_Pop_mioi_oswt_unreg;
  output dma_read_chnl_Pop_mioi_bawt;
  output dma_read_chnl_Pop_mioi_wen_comp;
  output [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt;
  input [63:0] dma_read_chnl_Pop_mioi_return_rsc_z;
  input dma_read_chnl_Pop_mioi_biwt;
  input dma_read_chnl_Pop_mioi_bdwt;


  // Interconnect Declarations
  reg dma_read_chnl_Pop_mioi_bcwt;
  reg [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_bfwt_31_0;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_chnl_Pop_mioi_bawt = dma_read_chnl_Pop_mioi_biwt | dma_read_chnl_Pop_mioi_bcwt;
  assign dma_read_chnl_Pop_mioi_wen_comp = (~ dma_read_chnl_Pop_mioi_oswt_unreg)
      | dma_read_chnl_Pop_mioi_bawt;
  assign dma_read_chnl_Pop_mioi_return_rsc_z_mxwt = MUX_v_32_2_2((dma_read_chnl_Pop_mioi_return_rsc_z[31:0]),
      dma_read_chnl_Pop_mioi_return_rsc_z_bfwt_31_0, dma_read_chnl_Pop_mioi_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_chnl_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_read_chnl_Pop_mioi_bcwt <= ~((~(dma_read_chnl_Pop_mioi_bcwt | dma_read_chnl_Pop_mioi_biwt))
          | dma_read_chnl_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( dma_read_chnl_Pop_mioi_biwt ) begin
      dma_read_chnl_Pop_mioi_return_rsc_z_bfwt_31_0 <= dma_read_chnl_Pop_mioi_return_rsc_z[31:0];
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl
    (
  clk, rst, load_wen, load_wten, dma_read_chnl_Pop_mioi_oswt_unreg, dma_read_chnl_Pop_mioi_iswt0,
      dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_psct, dma_read_chnl_Pop_mioi_biwt,
      dma_read_chnl_Pop_mioi_bdwt, dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_sct,
      dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld, dma_read_chnl_Pop_mioi_iswt0_pff
);
  input clk;
  input rst;
  input load_wen;
  input load_wten;
  input dma_read_chnl_Pop_mioi_oswt_unreg;
  input dma_read_chnl_Pop_mioi_iswt0;
  input dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_psct;
  output dma_read_chnl_Pop_mioi_biwt;
  output dma_read_chnl_Pop_mioi_bdwt;
  output dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_sct;
  input dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld;
  input dma_read_chnl_Pop_mioi_iswt0_pff;


  // Interconnect Declarations
  wire dma_read_chnl_Pop_mioi_ogwt;
  reg dma_read_chnl_Pop_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_chnl_Pop_mioi_bdwt = dma_read_chnl_Pop_mioi_oswt_unreg & load_wen;
  assign dma_read_chnl_Pop_mioi_biwt = dma_read_chnl_Pop_mioi_ogwt & dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld;
  assign dma_read_chnl_Pop_mioi_ogwt = ((~ load_wten) & dma_read_chnl_Pop_mioi_iswt0)
      | dma_read_chnl_Pop_mioi_icwt;
  assign dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_sct = dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_psct
      & load_wen & dma_read_chnl_Pop_mioi_iswt0_pff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_chnl_Pop_mioi_icwt <= 1'b0;
    end
    else begin
      dma_read_chnl_Pop_mioi_icwt <= dma_read_chnl_Pop_mioi_ogwt & (~ dma_read_chnl_Pop_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp
    (
  clk, rst, dma_read_ctrl_Push_mioi_oswt_unreg, dma_read_ctrl_Push_mioi_bawt, dma_read_ctrl_Push_mioi_wen_comp,
      dma_read_ctrl_Push_mioi_biwt, dma_read_ctrl_Push_mioi_bdwt
);
  input clk;
  input rst;
  input dma_read_ctrl_Push_mioi_oswt_unreg;
  output dma_read_ctrl_Push_mioi_bawt;
  output dma_read_ctrl_Push_mioi_wen_comp;
  input dma_read_ctrl_Push_mioi_biwt;
  input dma_read_ctrl_Push_mioi_bdwt;


  // Interconnect Declarations
  reg dma_read_ctrl_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_ctrl_Push_mioi_bawt = dma_read_ctrl_Push_mioi_biwt | dma_read_ctrl_Push_mioi_bcwt;
  assign dma_read_ctrl_Push_mioi_wen_comp = (~ dma_read_ctrl_Push_mioi_oswt_unreg)
      | dma_read_ctrl_Push_mioi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_read_ctrl_Push_mioi_bcwt <= ~((~(dma_read_ctrl_Push_mioi_bcwt | dma_read_ctrl_Push_mioi_biwt))
          | dma_read_ctrl_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl
    (
  clk, rst, load_wen, dma_read_ctrl_Push_mioi_oswt_unreg, dma_read_ctrl_Push_mioi_iswt0,
      load_wten, dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_psct, dma_read_ctrl_Push_mioi_biwt,
      dma_read_ctrl_Push_mioi_bdwt, dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_sct,
      dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld, dma_read_ctrl_Push_mioi_iswt0_pff
);
  input clk;
  input rst;
  input load_wen;
  input dma_read_ctrl_Push_mioi_oswt_unreg;
  input dma_read_ctrl_Push_mioi_iswt0;
  input load_wten;
  input dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_psct;
  output dma_read_ctrl_Push_mioi_biwt;
  output dma_read_ctrl_Push_mioi_bdwt;
  output dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_sct;
  input dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  input dma_read_ctrl_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire dma_read_ctrl_Push_mioi_ogwt;
  reg dma_read_ctrl_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_ctrl_Push_mioi_bdwt = dma_read_ctrl_Push_mioi_oswt_unreg & load_wen;
  assign dma_read_ctrl_Push_mioi_biwt = dma_read_ctrl_Push_mioi_ogwt & dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  assign dma_read_ctrl_Push_mioi_ogwt = ((~ load_wten) & dma_read_ctrl_Push_mioi_iswt0)
      | dma_read_ctrl_Push_mioi_icwt;
  assign dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_sct = dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_psct
      & load_wen & dma_read_ctrl_Push_mioi_iswt0_pff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_Push_mioi_icwt <= 1'b0;
    end
    else begin
      dma_read_ctrl_Push_mioi_icwt <= dma_read_ctrl_Push_mioi_ogwt & (~ dma_read_ctrl_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_config_config_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_config_config_fsm (
  clk, rst, fsm_output, CONFIG_LOOP_C_0_tr0
);
  input clk;
  input rst;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;
  input CONFIG_LOOP_C_0_tr0;


  // FSM State Type Declaration for esp_acc_softmax_sysc_softmax_sysc_config_config_fsm_1
  parameter
    config_rlp_C_0 = 2'd0,
    CONFIG_LOOP_C_0 = 2'd1,
    CONFIG_DONE_LOOP_C_0 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_softmax_sysc_softmax_sysc_config_config_fsm_1
    case (state_var)
      CONFIG_LOOP_C_0 : begin
        fsm_output = 3'b010;
        if ( CONFIG_LOOP_C_0_tr0 ) begin
          state_var_NS = CONFIG_LOOP_C_0;
        end
        else begin
          state_var_NS = CONFIG_DONE_LOOP_C_0;
        end
      end
      CONFIG_DONE_LOOP_C_0 : begin
        fsm_output = 3'b100;
        state_var_NS = CONFIG_DONE_LOOP_C_0;
      end
      // config_rlp_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = CONFIG_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= config_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_req_obj
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_req_obj (
  clk, rst, plm_out_cns_req_vz, store_wen, plm_out_cns_req_obj_oswt_unreg, plm_out_cns_req_obj_bawt,
      plm_out_cns_req_obj_iswt0, plm_out_cns_req_obj_wen_comp
);
  input clk;
  input rst;
  input plm_out_cns_req_vz;
  input store_wen;
  input plm_out_cns_req_obj_oswt_unreg;
  output plm_out_cns_req_obj_bawt;
  input plm_out_cns_req_obj_iswt0;
  output plm_out_cns_req_obj_wen_comp;


  // Interconnect Declarations
  wire plm_out_cns_req_obj_vd;
  wire plm_out_cns_req_obj_biwt;
  wire plm_out_cns_req_obj_bdwt;
  wire plm_out_cns_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_mgc_in_sync_v2 #(.valid(32'sd1)) plm_out_cns_req_obj (
      .vd(plm_out_cns_req_obj_vd),
      .vz(plm_out_cns_req_vz)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl
      softmax_sysc_store_store_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl_inst
      (
      .store_wen(store_wen),
      .plm_out_cns_req_obj_oswt_unreg(plm_out_cns_req_obj_oswt_unreg),
      .plm_out_cns_req_obj_iswt0(plm_out_cns_req_obj_iswt0),
      .plm_out_cns_req_obj_vd(plm_out_cns_req_obj_vd),
      .plm_out_cns_req_obj_biwt(plm_out_cns_req_obj_biwt),
      .plm_out_cns_req_obj_bdwt(plm_out_cns_req_obj_bdwt),
      .plm_out_cns_req_obj_bcwt(plm_out_cns_req_obj_bcwt)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_req_obj_plm_out_cns_req_wait_dp
      softmax_sysc_store_store_plm_out_cns_req_obj_plm_out_cns_req_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_req_obj_oswt_unreg(plm_out_cns_req_obj_oswt_unreg),
      .plm_out_cns_req_obj_bawt(plm_out_cns_req_obj_bawt),
      .plm_out_cns_req_obj_wen_comp(plm_out_cns_req_obj_wen_comp),
      .plm_out_cns_req_obj_biwt(plm_out_cns_req_obj_biwt),
      .plm_out_cns_req_obj_bdwt(plm_out_cns_req_obj_bdwt),
      .plm_out_cns_req_obj_bcwt(plm_out_cns_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_rls_obj
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_rls_obj (
  clk, rst, plm_out_cns_rls_lz, store_wen, store_wten, plm_out_cns_rls_obj_oswt_unreg,
      plm_out_cns_rls_obj_bawt, plm_out_cns_rls_obj_iswt0
);
  input clk;
  input rst;
  output plm_out_cns_rls_lz;
  input store_wen;
  input store_wten;
  input plm_out_cns_rls_obj_oswt_unreg;
  output plm_out_cns_rls_obj_bawt;
  input plm_out_cns_rls_obj_iswt0;


  // Interconnect Declarations
  wire plm_out_cns_rls_obj_biwt;
  wire plm_out_cns_rls_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_mgc_io_sync_v2 #(.valid(32'sd0)) plm_out_cns_rls_obj (
      .ld(plm_out_cns_rls_obj_biwt),
      .lz(plm_out_cns_rls_lz)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl
      softmax_sysc_store_store_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl_inst
      (
      .store_wen(store_wen),
      .store_wten(store_wten),
      .plm_out_cns_rls_obj_oswt_unreg(plm_out_cns_rls_obj_oswt_unreg),
      .plm_out_cns_rls_obj_iswt0(plm_out_cns_rls_obj_iswt0),
      .plm_out_cns_rls_obj_biwt(plm_out_cns_rls_obj_biwt),
      .plm_out_cns_rls_obj_bdwt(plm_out_cns_rls_obj_bdwt)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_rls_obj_plm_out_cns_rls_wait_dp
      softmax_sysc_store_store_plm_out_cns_rls_obj_plm_out_cns_rls_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_rls_obj_bawt(plm_out_cns_rls_obj_bawt),
      .plm_out_cns_rls_obj_biwt(plm_out_cns_rls_obj_biwt),
      .plm_out_cns_rls_obj_bdwt(plm_out_cns_rls_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cnsi_1
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cnsi_1 (
  clk, rst, plm_out_cnsi_q_d, plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d, store_wen,
      store_wten, plm_out_cnsi_oswt_unreg, plm_out_cnsi_bawt, plm_out_cnsi_iswt0,
      plm_out_cnsi_q_d_mxwt, plm_out_cnsi_iswt0_pff
);
  input clk;
  input rst;
  input [31:0] plm_out_cnsi_q_d;
  output plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d;
  input store_wen;
  input store_wten;
  input plm_out_cnsi_oswt_unreg;
  output plm_out_cnsi_bawt;
  input plm_out_cnsi_iswt0;
  output [31:0] plm_out_cnsi_q_d_mxwt;
  input plm_out_cnsi_iswt0_pff;


  // Interconnect Declarations
  wire plm_out_cnsi_biwt;
  wire plm_out_cnsi_bdwt;
  wire plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_store_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cnsi_1_plm_out_cns_wait_ctrl
      softmax_sysc_store_store_plm_out_cnsi_1_plm_out_cns_wait_ctrl_inst (
      .store_wen(store_wen),
      .store_wten(store_wten),
      .plm_out_cnsi_oswt_unreg(plm_out_cnsi_oswt_unreg),
      .plm_out_cnsi_iswt0(plm_out_cnsi_iswt0),
      .plm_out_cnsi_biwt(plm_out_cnsi_biwt),
      .plm_out_cnsi_bdwt(plm_out_cnsi_bdwt),
      .plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_store_sct(plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_store_sct),
      .plm_out_cnsi_iswt0_pff(plm_out_cnsi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cnsi_1_plm_out_cns_wait_dp
      softmax_sysc_store_store_plm_out_cnsi_1_plm_out_cns_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_out_cnsi_q_d(plm_out_cnsi_q_d),
      .plm_out_cnsi_bawt(plm_out_cnsi_bawt),
      .plm_out_cnsi_q_d_mxwt(plm_out_cnsi_q_d_mxwt),
      .plm_out_cnsi_biwt(plm_out_cnsi_biwt),
      .plm_out_cnsi_bdwt(plm_out_cnsi_bdwt)
    );
  assign plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d = plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_store_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_chnl_Push_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_chnl_Push_mioi (
  clk, rst, dma_write_chnl_val, dma_write_chnl_rdy, dma_write_chnl_msg, store_wen,
      store_wten, dma_write_chnl_Push_mioi_m_rsc_dat, dma_write_chnl_Push_mioi_oswt_unreg,
      dma_write_chnl_Push_mioi_bawt, dma_write_chnl_Push_mioi_iswt0, dma_write_chnl_Push_mioi_wen_comp,
      dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct, dma_write_chnl_Push_mioi_iswt0_pff
);
  input clk;
  input rst;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;
  input store_wen;
  input store_wten;
  input [63:0] dma_write_chnl_Push_mioi_m_rsc_dat;
  input dma_write_chnl_Push_mioi_oswt_unreg;
  output dma_write_chnl_Push_mioi_bawt;
  input dma_write_chnl_Push_mioi_iswt0;
  output dma_write_chnl_Push_mioi_wen_comp;
  input dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct;
  input dma_write_chnl_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire dma_write_chnl_Push_mioi_biwt;
  wire dma_write_chnl_Push_mioi_bdwt;
  wire dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_sct;
  wire dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  wire [63:0] nl_dma_write_chnl_Push_mioi_m_rsc_dat;
  assign nl_dma_write_chnl_Push_mioi_m_rsc_dat = {32'b11011110101011011011111011101111
      , (dma_write_chnl_Push_mioi_m_rsc_dat[31:0])};
  esp_acc_softmax_sysc_Connections_OutBlocking_dma_data_t_Connections_SYN_PORT_Push
      dma_write_chnl_Push_mioi (
      .this_val(dma_write_chnl_val),
      .this_rdy(dma_write_chnl_rdy),
      .this_msg(dma_write_chnl_msg),
      .m_rsc_dat(nl_dma_write_chnl_Push_mioi_m_rsc_dat[63:0]),
      .ccs_ccore_start_rsc_dat(dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_sct),
      .ccs_ccore_done_sync_vld(dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl
      softmax_sysc_store_store_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .store_wen(store_wen),
      .store_wten(store_wten),
      .dma_write_chnl_Push_mioi_oswt_unreg(dma_write_chnl_Push_mioi_oswt_unreg),
      .dma_write_chnl_Push_mioi_iswt0(dma_write_chnl_Push_mioi_iswt0),
      .dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct(dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct),
      .dma_write_chnl_Push_mioi_biwt(dma_write_chnl_Push_mioi_biwt),
      .dma_write_chnl_Push_mioi_bdwt(dma_write_chnl_Push_mioi_bdwt),
      .dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_sct(dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_sct),
      .dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld(dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld),
      .dma_write_chnl_Push_mioi_iswt0_pff(dma_write_chnl_Push_mioi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp
      softmax_sysc_store_store_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_chnl_Push_mioi_oswt_unreg(dma_write_chnl_Push_mioi_oswt_unreg),
      .dma_write_chnl_Push_mioi_bawt(dma_write_chnl_Push_mioi_bawt),
      .dma_write_chnl_Push_mioi_wen_comp(dma_write_chnl_Push_mioi_wen_comp),
      .dma_write_chnl_Push_mioi_biwt(dma_write_chnl_Push_mioi_biwt),
      .dma_write_chnl_Push_mioi_bdwt(dma_write_chnl_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_ctrl_Push_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_ctrl_Push_mioi (
  clk, rst, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg, store_wen,
      store_wten, dma_write_ctrl_Push_mioi_m_index_rsc_dat, dma_write_ctrl_Push_mioi_oswt_unreg,
      dma_write_ctrl_Push_mioi_bawt, dma_write_ctrl_Push_mioi_iswt0, dma_write_ctrl_Push_mioi_wen_comp,
      dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct, dma_write_ctrl_Push_mioi_iswt0_pff
);
  input clk;
  input rst;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  input store_wen;
  input store_wten;
  input [31:0] dma_write_ctrl_Push_mioi_m_index_rsc_dat;
  input dma_write_ctrl_Push_mioi_oswt_unreg;
  output dma_write_ctrl_Push_mioi_bawt;
  input dma_write_ctrl_Push_mioi_iswt0;
  output dma_write_ctrl_Push_mioi_wen_comp;
  input dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct;
  input dma_write_ctrl_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire dma_write_ctrl_Push_mioi_biwt;
  wire dma_write_ctrl_Push_mioi_bdwt;
  wire dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_sct;
  wire dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_dma_write_ctrl_Push_mioi_m_index_rsc_dat;
  assign nl_dma_write_ctrl_Push_mioi_m_index_rsc_dat = {(dma_write_ctrl_Push_mioi_m_index_rsc_dat[31:7])
      , 7'b0000000};
  esp_acc_softmax_sysc_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push
      dma_write_ctrl_Push_mioi (
      .this_val(dma_write_ctrl_val),
      .this_rdy(dma_write_ctrl_rdy),
      .this_msg(dma_write_ctrl_msg),
      .m_index_rsc_dat(nl_dma_write_ctrl_Push_mioi_m_index_rsc_dat[31:0]),
      .ccs_ccore_start_rsc_dat(dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_sct),
      .ccs_ccore_done_sync_vld(dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl
      softmax_sysc_store_store_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .store_wen(store_wen),
      .store_wten(store_wten),
      .dma_write_ctrl_Push_mioi_oswt_unreg(dma_write_ctrl_Push_mioi_oswt_unreg),
      .dma_write_ctrl_Push_mioi_iswt0(dma_write_ctrl_Push_mioi_iswt0),
      .dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct(dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct),
      .dma_write_ctrl_Push_mioi_biwt(dma_write_ctrl_Push_mioi_biwt),
      .dma_write_ctrl_Push_mioi_bdwt(dma_write_ctrl_Push_mioi_bdwt),
      .dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_sct(dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_sct),
      .dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld(dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .dma_write_ctrl_Push_mioi_iswt0_pff(dma_write_ctrl_Push_mioi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp
      softmax_sysc_store_store_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_ctrl_Push_mioi_oswt_unreg(dma_write_ctrl_Push_mioi_oswt_unreg),
      .dma_write_ctrl_Push_mioi_bawt(dma_write_ctrl_Push_mioi_bawt),
      .dma_write_ctrl_Push_mioi_wen_comp(dma_write_ctrl_Push_mioi_wen_comp),
      .dma_write_ctrl_Push_mioi_biwt(dma_write_ctrl_Push_mioi_biwt),
      .dma_write_ctrl_Push_mioi_bdwt(dma_write_ctrl_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store_output_ready_ack_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store_output_ready_ack_mioi (
  clk, rst, output_ready_req_req, output_ready_ack_ack, store_wen, output_ready_ack_mioi_oswt_unreg,
      output_ready_ack_mioi_bawt, output_ready_ack_mioi_iswt0, store_wten, output_ready_ack_mioi_wen_comp,
      output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_psct, output_ready_ack_mioi_iswt0_pff
);
  input clk;
  input rst;
  input output_ready_req_req;
  output output_ready_ack_ack;
  input store_wen;
  input output_ready_ack_mioi_oswt_unreg;
  output output_ready_ack_mioi_bawt;
  input output_ready_ack_mioi_iswt0;
  input store_wten;
  output output_ready_ack_mioi_wen_comp;
  input output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_psct;
  input output_ready_ack_mioi_iswt0_pff;


  // Interconnect Declarations
  wire output_ready_ack_mioi_biwt;
  wire output_ready_ack_mioi_bdwt;
  wire output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_sct;
  wire output_ready_ack_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_handshake_t_ack  output_ready_ack_mioi (
      .this_req_req(output_ready_req_req),
      .this_ack_ack(output_ready_ack_ack),
      .ccs_ccore_start_rsc_dat(output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_sct),
      .ccs_ccore_done_sync_vld(output_ready_ack_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_output_ready_ack_mioi_output_ready_ack_mio_wait_ctrl
      softmax_sysc_store_store_output_ready_ack_mioi_output_ready_ack_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .store_wen(store_wen),
      .output_ready_ack_mioi_oswt_unreg(output_ready_ack_mioi_oswt_unreg),
      .output_ready_ack_mioi_iswt0(output_ready_ack_mioi_iswt0),
      .store_wten(store_wten),
      .output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_psct(output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_psct),
      .output_ready_ack_mioi_biwt(output_ready_ack_mioi_biwt),
      .output_ready_ack_mioi_bdwt(output_ready_ack_mioi_bdwt),
      .output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_sct(output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_sct),
      .output_ready_ack_mioi_ccs_ccore_done_sync_vld(output_ready_ack_mioi_ccs_ccore_done_sync_vld),
      .output_ready_ack_mioi_iswt0_pff(output_ready_ack_mioi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_output_ready_ack_mioi_output_ready_ack_mio_wait_dp
      softmax_sysc_store_store_output_ready_ack_mioi_output_ready_ack_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .output_ready_ack_mioi_oswt_unreg(output_ready_ack_mioi_oswt_unreg),
      .output_ready_ack_mioi_bawt(output_ready_ack_mioi_bawt),
      .output_ready_ack_mioi_wen_comp(output_ready_ack_mioi_wen_comp),
      .output_ready_ack_mioi_biwt(output_ready_ack_mioi_biwt),
      .output_ready_ack_mioi_bdwt(output_ready_ack_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_req_obj
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_req_obj (
  clk, rst, plm_out_cns_req_vz, compute_wen, plm_out_cns_req_obj_oswt_unreg, plm_out_cns_req_obj_bawt,
      plm_out_cns_req_obj_iswt0, plm_out_cns_req_obj_wen_comp
);
  input clk;
  input rst;
  input plm_out_cns_req_vz;
  input compute_wen;
  input plm_out_cns_req_obj_oswt_unreg;
  output plm_out_cns_req_obj_bawt;
  input plm_out_cns_req_obj_iswt0;
  output plm_out_cns_req_obj_wen_comp;


  // Interconnect Declarations
  wire plm_out_cns_req_obj_vd;
  wire plm_out_cns_req_obj_biwt;
  wire plm_out_cns_req_obj_bdwt;
  wire plm_out_cns_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_mgc_in_sync_v2 #(.valid(32'sd1)) plm_out_cns_req_obj (
      .vd(plm_out_cns_req_obj_vd),
      .vz(plm_out_cns_req_vz)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl
      softmax_sysc_compute_compute_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl_inst
      (
      .compute_wen(compute_wen),
      .plm_out_cns_req_obj_oswt_unreg(plm_out_cns_req_obj_oswt_unreg),
      .plm_out_cns_req_obj_iswt0(plm_out_cns_req_obj_iswt0),
      .plm_out_cns_req_obj_vd(plm_out_cns_req_obj_vd),
      .plm_out_cns_req_obj_biwt(plm_out_cns_req_obj_biwt),
      .plm_out_cns_req_obj_bdwt(plm_out_cns_req_obj_bdwt),
      .plm_out_cns_req_obj_bcwt(plm_out_cns_req_obj_bcwt)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_req_obj_plm_out_cns_req_wait_dp
      softmax_sysc_compute_compute_plm_out_cns_req_obj_plm_out_cns_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_req_obj_oswt_unreg(plm_out_cns_req_obj_oswt_unreg),
      .plm_out_cns_req_obj_bawt(plm_out_cns_req_obj_bawt),
      .plm_out_cns_req_obj_wen_comp(plm_out_cns_req_obj_wen_comp),
      .plm_out_cns_req_obj_biwt(plm_out_cns_req_obj_biwt),
      .plm_out_cns_req_obj_bdwt(plm_out_cns_req_obj_bdwt),
      .plm_out_cns_req_obj_bcwt(plm_out_cns_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_req_obj
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_req_obj (
  clk, rst, plm_in_cns_req_vz, compute_wen, plm_in_cns_req_obj_oswt_unreg, plm_in_cns_req_obj_bawt,
      plm_in_cns_req_obj_iswt0, plm_in_cns_req_obj_wen_comp
);
  input clk;
  input rst;
  input plm_in_cns_req_vz;
  input compute_wen;
  input plm_in_cns_req_obj_oswt_unreg;
  output plm_in_cns_req_obj_bawt;
  input plm_in_cns_req_obj_iswt0;
  output plm_in_cns_req_obj_wen_comp;


  // Interconnect Declarations
  wire plm_in_cns_req_obj_vd;
  wire plm_in_cns_req_obj_biwt;
  wire plm_in_cns_req_obj_bdwt;
  wire plm_in_cns_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_mgc_in_sync_v2 #(.valid(32'sd1)) plm_in_cns_req_obj (
      .vd(plm_in_cns_req_obj_vd),
      .vz(plm_in_cns_req_vz)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl
      softmax_sysc_compute_compute_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl_inst
      (
      .compute_wen(compute_wen),
      .plm_in_cns_req_obj_oswt_unreg(plm_in_cns_req_obj_oswt_unreg),
      .plm_in_cns_req_obj_iswt0(plm_in_cns_req_obj_iswt0),
      .plm_in_cns_req_obj_vd(plm_in_cns_req_obj_vd),
      .plm_in_cns_req_obj_biwt(plm_in_cns_req_obj_biwt),
      .plm_in_cns_req_obj_bdwt(plm_in_cns_req_obj_bdwt),
      .plm_in_cns_req_obj_bcwt(plm_in_cns_req_obj_bcwt)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_req_obj_plm_in_cns_req_wait_dp
      softmax_sysc_compute_compute_plm_in_cns_req_obj_plm_in_cns_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_req_obj_oswt_unreg(plm_in_cns_req_obj_oswt_unreg),
      .plm_in_cns_req_obj_bawt(plm_in_cns_req_obj_bawt),
      .plm_in_cns_req_obj_wen_comp(plm_in_cns_req_obj_wen_comp),
      .plm_in_cns_req_obj_biwt(plm_in_cns_req_obj_biwt),
      .plm_in_cns_req_obj_bdwt(plm_in_cns_req_obj_bdwt),
      .plm_in_cns_req_obj_bcwt(plm_in_cns_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_rls_obj
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_rls_obj (
  clk, rst, plm_in_cns_rls_lz, compute_wen, compute_wten, plm_in_cns_rls_obj_oswt_unreg,
      plm_in_cns_rls_obj_bawt, plm_in_cns_rls_obj_iswt0
);
  input clk;
  input rst;
  output plm_in_cns_rls_lz;
  input compute_wen;
  input compute_wten;
  input plm_in_cns_rls_obj_oswt_unreg;
  output plm_in_cns_rls_obj_bawt;
  input plm_in_cns_rls_obj_iswt0;


  // Interconnect Declarations
  wire plm_in_cns_rls_obj_biwt;
  wire plm_in_cns_rls_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_mgc_io_sync_v2 #(.valid(32'sd0)) plm_in_cns_rls_obj (
      .ld(plm_in_cns_rls_obj_biwt),
      .lz(plm_in_cns_rls_lz)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl
      softmax_sysc_compute_compute_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl_inst
      (
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .plm_in_cns_rls_obj_oswt_unreg(plm_in_cns_rls_obj_oswt_unreg),
      .plm_in_cns_rls_obj_iswt0(plm_in_cns_rls_obj_iswt0),
      .plm_in_cns_rls_obj_biwt(plm_in_cns_rls_obj_biwt),
      .plm_in_cns_rls_obj_bdwt(plm_in_cns_rls_obj_bdwt)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_rls_obj_plm_in_cns_rls_wait_dp
      softmax_sysc_compute_compute_plm_in_cns_rls_obj_plm_in_cns_rls_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_rls_obj_bawt(plm_in_cns_rls_obj_bawt),
      .plm_in_cns_rls_obj_biwt(plm_in_cns_rls_obj_biwt),
      .plm_in_cns_rls_obj_bdwt(plm_in_cns_rls_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp
    (
  clk, rst, compute_wen, compute_wten, CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg, CALC_SOFTMAX_LOOP_mul_cmp_bawt,
      CALC_SOFTMAX_LOOP_mul_cmp_iswt2, CALC_SOFTMAX_LOOP_mul_cmp_a_compute, CALC_SOFTMAX_LOOP_mul_cmp_b_compute,
      CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt
);
  input clk;
  input rst;
  input compute_wen;
  input compute_wten;
  input CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg;
  output CALC_SOFTMAX_LOOP_mul_cmp_bawt;
  input CALC_SOFTMAX_LOOP_mul_cmp_iswt2;
  input [66:0] CALC_SOFTMAX_LOOP_mul_cmp_a_compute;
  input [93:0] CALC_SOFTMAX_LOOP_mul_cmp_b_compute;
  output [31:0] CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt;


  // Interconnect Declarations
  wire CALC_SOFTMAX_LOOP_mul_cmp_biwt;
  wire CALC_SOFTMAX_LOOP_mul_cmp_bdwt;
  wire [94:0] CALC_SOFTMAX_LOOP_mul_cmp_z;
  wire [31:0] CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_mgc_mul_pipe #(.width_a(32'sd67),
  .signd_a(32'sd0),
  .width_b(32'sd94),
  .signd_b(32'sd0),
  .width_z(32'sd95),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) CALC_SOFTMAX_LOOP_mul_cmp (
      .a(CALC_SOFTMAX_LOOP_mul_cmp_a_compute),
      .b(CALC_SOFTMAX_LOOP_mul_cmp_b_compute),
      .clk(clk),
      .en(1'b1),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(CALC_SOFTMAX_LOOP_mul_cmp_z)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_ctrl
      softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg(CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg),
      .CALC_SOFTMAX_LOOP_mul_cmp_iswt2(CALC_SOFTMAX_LOOP_mul_cmp_iswt2),
      .CALC_SOFTMAX_LOOP_mul_cmp_biwt(CALC_SOFTMAX_LOOP_mul_cmp_biwt),
      .CALC_SOFTMAX_LOOP_mul_cmp_bdwt(CALC_SOFTMAX_LOOP_mul_cmp_bdwt)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_dp
      softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .CALC_SOFTMAX_LOOP_mul_cmp_bawt(CALC_SOFTMAX_LOOP_mul_cmp_bawt),
      .CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt(CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt_pconst),
      .CALC_SOFTMAX_LOOP_mul_cmp_biwt(CALC_SOFTMAX_LOOP_mul_cmp_biwt),
      .CALC_SOFTMAX_LOOP_mul_cmp_bdwt(CALC_SOFTMAX_LOOP_mul_cmp_bdwt),
      .CALC_SOFTMAX_LOOP_mul_cmp_z(CALC_SOFTMAX_LOOP_mul_cmp_z)
    );
  assign CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt = CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_rls_obj
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_rls_obj (
  clk, rst, plm_out_cns_rls_lz, compute_wen, compute_wten, plm_out_cns_rls_obj_oswt_unreg,
      plm_out_cns_rls_obj_bawt, plm_out_cns_rls_obj_iswt0
);
  input clk;
  input rst;
  output plm_out_cns_rls_lz;
  input compute_wen;
  input compute_wten;
  input plm_out_cns_rls_obj_oswt_unreg;
  output plm_out_cns_rls_obj_bawt;
  input plm_out_cns_rls_obj_iswt0;


  // Interconnect Declarations
  wire plm_out_cns_rls_obj_biwt;
  wire plm_out_cns_rls_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_mgc_io_sync_v2 #(.valid(32'sd0)) plm_out_cns_rls_obj (
      .ld(plm_out_cns_rls_obj_biwt),
      .lz(plm_out_cns_rls_lz)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl
      softmax_sysc_compute_compute_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl_inst
      (
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .plm_out_cns_rls_obj_oswt_unreg(plm_out_cns_rls_obj_oswt_unreg),
      .plm_out_cns_rls_obj_iswt0(plm_out_cns_rls_obj_iswt0),
      .plm_out_cns_rls_obj_biwt(plm_out_cns_rls_obj_biwt),
      .plm_out_cns_rls_obj_bdwt(plm_out_cns_rls_obj_bdwt)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_rls_obj_plm_out_cns_rls_wait_dp
      softmax_sysc_compute_compute_plm_out_cns_rls_obj_plm_out_cns_rls_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_rls_obj_bawt(plm_out_cns_rls_obj_bawt),
      .plm_out_cns_rls_obj_biwt(plm_out_cns_rls_obj_biwt),
      .plm_out_cns_rls_obj_bdwt(plm_out_cns_rls_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cnsi_1
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cnsi_1 (
  clk, rst, compute_wen, compute_wten, plm_out_cnsi_oswt_unreg, plm_out_cnsi_bawt,
      plm_out_cnsi_iswt0, plm_out_cnsi_we_d_pff, plm_out_cnsi_iswt0_pff
);
  input clk;
  input rst;
  input compute_wen;
  input compute_wten;
  input plm_out_cnsi_oswt_unreg;
  output plm_out_cnsi_bawt;
  input plm_out_cnsi_iswt0;
  output plm_out_cnsi_we_d_pff;
  input plm_out_cnsi_iswt0_pff;


  // Interconnect Declarations
  wire plm_out_cnsi_biwt;
  wire plm_out_cnsi_bdwt;
  wire plm_out_cnsi_we_d_compute_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cnsi_1_plm_out_cns_wait_ctrl
      softmax_sysc_compute_compute_plm_out_cnsi_1_plm_out_cns_wait_ctrl_inst (
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .plm_out_cnsi_oswt_unreg(plm_out_cnsi_oswt_unreg),
      .plm_out_cnsi_iswt0(plm_out_cnsi_iswt0),
      .plm_out_cnsi_biwt(plm_out_cnsi_biwt),
      .plm_out_cnsi_bdwt(plm_out_cnsi_bdwt),
      .plm_out_cnsi_we_d_compute_sct_pff(plm_out_cnsi_we_d_compute_sct_iff),
      .plm_out_cnsi_iswt0_pff(plm_out_cnsi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cnsi_1_plm_out_cns_wait_dp
      softmax_sysc_compute_compute_plm_out_cnsi_1_plm_out_cns_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_out_cnsi_bawt(plm_out_cnsi_bawt),
      .plm_out_cnsi_biwt(plm_out_cnsi_biwt),
      .plm_out_cnsi_bdwt(plm_out_cnsi_bdwt)
    );
  assign plm_out_cnsi_we_d_pff = plm_out_cnsi_we_d_compute_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cnsi_1
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cnsi_1 (
  clk, rst, plm_in_cnsi_q_d, plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d, compute_wen,
      compute_wten, plm_in_cnsi_oswt_unreg, plm_in_cnsi_bawt, plm_in_cnsi_iswt0,
      plm_in_cnsi_q_d_mxwt, plm_in_cnsi_iswt0_pff
);
  input clk;
  input rst;
  input [31:0] plm_in_cnsi_q_d;
  output plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d;
  input compute_wen;
  input compute_wten;
  input plm_in_cnsi_oswt_unreg;
  output plm_in_cnsi_bawt;
  input plm_in_cnsi_iswt0;
  output [31:0] plm_in_cnsi_q_d_mxwt;
  input plm_in_cnsi_iswt0_pff;


  // Interconnect Declarations
  wire plm_in_cnsi_biwt;
  wire plm_in_cnsi_bdwt;
  wire plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_compute_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cnsi_1_plm_in_cns_wait_ctrl
      softmax_sysc_compute_compute_plm_in_cnsi_1_plm_in_cns_wait_ctrl_inst (
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .plm_in_cnsi_oswt_unreg(plm_in_cnsi_oswt_unreg),
      .plm_in_cnsi_iswt0(plm_in_cnsi_iswt0),
      .plm_in_cnsi_biwt(plm_in_cnsi_biwt),
      .plm_in_cnsi_bdwt(plm_in_cnsi_bdwt),
      .plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_compute_sct(plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_compute_sct),
      .plm_in_cnsi_iswt0_pff(plm_in_cnsi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cnsi_1_plm_in_cns_wait_dp
      softmax_sysc_compute_compute_plm_in_cnsi_1_plm_in_cns_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_in_cnsi_q_d(plm_in_cnsi_q_d),
      .plm_in_cnsi_bawt(plm_in_cnsi_bawt),
      .plm_in_cnsi_q_d_mxwt(plm_in_cnsi_q_d_mxwt),
      .plm_in_cnsi_biwt(plm_in_cnsi_biwt),
      .plm_in_cnsi_bdwt(plm_in_cnsi_bdwt)
    );
  assign plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d = plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_compute_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_output_ready_req_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_output_ready_req_mioi (
  clk, rst, output_ready_req_req, output_ready_ack_ack, compute_wen, compute_wten,
      output_ready_req_mioi_oswt_unreg, output_ready_req_mioi_bawt, output_ready_req_mioi_iswt0,
      output_ready_req_mioi_wen_comp, output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_psct,
      output_ready_req_mioi_iswt0_pff
);
  input clk;
  input rst;
  output output_ready_req_req;
  input output_ready_ack_ack;
  input compute_wen;
  input compute_wten;
  input output_ready_req_mioi_oswt_unreg;
  output output_ready_req_mioi_bawt;
  input output_ready_req_mioi_iswt0;
  output output_ready_req_mioi_wen_comp;
  input output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_psct;
  input output_ready_req_mioi_iswt0_pff;


  // Interconnect Declarations
  wire output_ready_req_mioi_biwt;
  wire output_ready_req_mioi_bdwt;
  wire output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_sct;
  wire output_ready_req_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_handshake_t_req  output_ready_req_mioi (
      .this_req_req(output_ready_req_req),
      .this_ack_ack(output_ready_ack_ack),
      .ccs_ccore_start_rsc_dat(output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_sct),
      .ccs_ccore_done_sync_vld(output_ready_req_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_output_ready_req_mioi_output_ready_req_mio_wait_ctrl
      softmax_sysc_compute_compute_output_ready_req_mioi_output_ready_req_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .output_ready_req_mioi_oswt_unreg(output_ready_req_mioi_oswt_unreg),
      .output_ready_req_mioi_iswt0(output_ready_req_mioi_iswt0),
      .output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_psct(output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_psct),
      .output_ready_req_mioi_biwt(output_ready_req_mioi_biwt),
      .output_ready_req_mioi_bdwt(output_ready_req_mioi_bdwt),
      .output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_sct(output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_sct),
      .output_ready_req_mioi_ccs_ccore_done_sync_vld(output_ready_req_mioi_ccs_ccore_done_sync_vld),
      .output_ready_req_mioi_iswt0_pff(output_ready_req_mioi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_output_ready_req_mioi_output_ready_req_mio_wait_dp
      softmax_sysc_compute_compute_output_ready_req_mioi_output_ready_req_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .output_ready_req_mioi_oswt_unreg(output_ready_req_mioi_oswt_unreg),
      .output_ready_req_mioi_bawt(output_ready_req_mioi_bawt),
      .output_ready_req_mioi_wen_comp(output_ready_req_mioi_wen_comp),
      .output_ready_req_mioi_biwt(output_ready_req_mioi_biwt),
      .output_ready_req_mioi_bdwt(output_ready_req_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_input_ready_ack_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_input_ready_ack_mioi (
  clk, rst, input_ready_req_req, input_ready_ack_ack, compute_wen, compute_wten,
      input_ready_ack_mioi_oswt_unreg, input_ready_ack_mioi_bawt, input_ready_ack_mioi_iswt0,
      input_ready_ack_mioi_wen_comp, input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_psct,
      input_ready_ack_mioi_iswt0_pff
);
  input clk;
  input rst;
  input input_ready_req_req;
  output input_ready_ack_ack;
  input compute_wen;
  input compute_wten;
  input input_ready_ack_mioi_oswt_unreg;
  output input_ready_ack_mioi_bawt;
  input input_ready_ack_mioi_iswt0;
  output input_ready_ack_mioi_wen_comp;
  input input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_psct;
  input input_ready_ack_mioi_iswt0_pff;


  // Interconnect Declarations
  wire input_ready_ack_mioi_biwt;
  wire input_ready_ack_mioi_bdwt;
  wire input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_sct;
  wire input_ready_ack_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_handshake_t_ack  input_ready_ack_mioi (
      .this_req_req(input_ready_req_req),
      .this_ack_ack(input_ready_ack_ack),
      .ccs_ccore_start_rsc_dat(input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_sct),
      .ccs_ccore_done_sync_vld(input_ready_ack_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_input_ready_ack_mioi_input_ready_ack_mio_wait_ctrl
      softmax_sysc_compute_compute_input_ready_ack_mioi_input_ready_ack_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .input_ready_ack_mioi_oswt_unreg(input_ready_ack_mioi_oswt_unreg),
      .input_ready_ack_mioi_iswt0(input_ready_ack_mioi_iswt0),
      .input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_psct(input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_psct),
      .input_ready_ack_mioi_biwt(input_ready_ack_mioi_biwt),
      .input_ready_ack_mioi_bdwt(input_ready_ack_mioi_bdwt),
      .input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_sct(input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_sct),
      .input_ready_ack_mioi_ccs_ccore_done_sync_vld(input_ready_ack_mioi_ccs_ccore_done_sync_vld),
      .input_ready_ack_mioi_iswt0_pff(input_ready_ack_mioi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_input_ready_ack_mioi_input_ready_ack_mio_wait_dp
      softmax_sysc_compute_compute_input_ready_ack_mioi_input_ready_ack_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_ready_ack_mioi_oswt_unreg(input_ready_ack_mioi_oswt_unreg),
      .input_ready_ack_mioi_bawt(input_ready_ack_mioi_bawt),
      .input_ready_ack_mioi_wen_comp(input_ready_ack_mioi_wen_comp),
      .input_ready_ack_mioi_biwt(input_ready_ack_mioi_biwt),
      .input_ready_ack_mioi_bdwt(input_ready_ack_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1
    (
  clk, rst, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      compute_wen, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0,
      compute_wten, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff
);
  input clk;
  input rst;
  input [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  input compute_wen;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0;
  input compute_wten;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1;
  output [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff;


  // Interconnect Declarations
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_compute_sct;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_compute_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_ctrl
      softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_ctrl_inst
      (
      .compute_wen(compute_wen),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0),
      .compute_wten(compute_wten),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_compute_sct(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_compute_sct),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_compute_sct_pff(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_compute_sct_iff),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_dp
      softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2)
    );
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_compute_sct_iff;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_compute_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_req_obj
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_req_obj (
  clk, rst, plm_in_cns_req_vz, load_wen, plm_in_cns_req_obj_oswt_unreg, plm_in_cns_req_obj_bawt,
      plm_in_cns_req_obj_iswt0, plm_in_cns_req_obj_wen_comp
);
  input clk;
  input rst;
  input plm_in_cns_req_vz;
  input load_wen;
  input plm_in_cns_req_obj_oswt_unreg;
  output plm_in_cns_req_obj_bawt;
  input plm_in_cns_req_obj_iswt0;
  output plm_in_cns_req_obj_wen_comp;


  // Interconnect Declarations
  wire plm_in_cns_req_obj_vd;
  wire plm_in_cns_req_obj_biwt;
  wire plm_in_cns_req_obj_bdwt;
  wire plm_in_cns_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_mgc_in_sync_v2 #(.valid(32'sd1)) plm_in_cns_req_obj (
      .vd(plm_in_cns_req_obj_vd),
      .vz(plm_in_cns_req_vz)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl
      softmax_sysc_load_load_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl_inst (
      .load_wen(load_wen),
      .plm_in_cns_req_obj_oswt_unreg(plm_in_cns_req_obj_oswt_unreg),
      .plm_in_cns_req_obj_iswt0(plm_in_cns_req_obj_iswt0),
      .plm_in_cns_req_obj_vd(plm_in_cns_req_obj_vd),
      .plm_in_cns_req_obj_biwt(plm_in_cns_req_obj_biwt),
      .plm_in_cns_req_obj_bdwt(plm_in_cns_req_obj_bdwt),
      .plm_in_cns_req_obj_bcwt(plm_in_cns_req_obj_bcwt)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_req_obj_plm_in_cns_req_wait_dp
      softmax_sysc_load_load_plm_in_cns_req_obj_plm_in_cns_req_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_req_obj_oswt_unreg(plm_in_cns_req_obj_oswt_unreg),
      .plm_in_cns_req_obj_bawt(plm_in_cns_req_obj_bawt),
      .plm_in_cns_req_obj_wen_comp(plm_in_cns_req_obj_wen_comp),
      .plm_in_cns_req_obj_biwt(plm_in_cns_req_obj_biwt),
      .plm_in_cns_req_obj_bdwt(plm_in_cns_req_obj_bdwt),
      .plm_in_cns_req_obj_bcwt(plm_in_cns_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_rls_obj
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_rls_obj (
  clk, rst, plm_in_cns_rls_lz, load_wen, load_wten, plm_in_cns_rls_obj_oswt_unreg,
      plm_in_cns_rls_obj_bawt, plm_in_cns_rls_obj_iswt0
);
  input clk;
  input rst;
  output plm_in_cns_rls_lz;
  input load_wen;
  input load_wten;
  input plm_in_cns_rls_obj_oswt_unreg;
  output plm_in_cns_rls_obj_bawt;
  input plm_in_cns_rls_obj_iswt0;


  // Interconnect Declarations
  wire plm_in_cns_rls_obj_biwt;
  wire plm_in_cns_rls_obj_bdwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_mgc_io_sync_v2 #(.valid(32'sd0)) plm_in_cns_rls_obj (
      .ld(plm_in_cns_rls_obj_biwt),
      .lz(plm_in_cns_rls_lz)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl
      softmax_sysc_load_load_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl_inst (
      .load_wen(load_wen),
      .load_wten(load_wten),
      .plm_in_cns_rls_obj_oswt_unreg(plm_in_cns_rls_obj_oswt_unreg),
      .plm_in_cns_rls_obj_iswt0(plm_in_cns_rls_obj_iswt0),
      .plm_in_cns_rls_obj_biwt(plm_in_cns_rls_obj_biwt),
      .plm_in_cns_rls_obj_bdwt(plm_in_cns_rls_obj_bdwt)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_rls_obj_plm_in_cns_rls_wait_dp
      softmax_sysc_load_load_plm_in_cns_rls_obj_plm_in_cns_rls_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_rls_obj_bawt(plm_in_cns_rls_obj_bawt),
      .plm_in_cns_rls_obj_biwt(plm_in_cns_rls_obj_biwt),
      .plm_in_cns_rls_obj_bdwt(plm_in_cns_rls_obj_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cnsi_1
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cnsi_1 (
  clk, rst, load_wen, load_wten, plm_in_cnsi_oswt_unreg, plm_in_cnsi_bawt, plm_in_cnsi_iswt0,
      plm_in_cnsi_we_d_pff, plm_in_cnsi_iswt0_pff
);
  input clk;
  input rst;
  input load_wen;
  input load_wten;
  input plm_in_cnsi_oswt_unreg;
  output plm_in_cnsi_bawt;
  input plm_in_cnsi_iswt0;
  output plm_in_cnsi_we_d_pff;
  input plm_in_cnsi_iswt0_pff;


  // Interconnect Declarations
  wire plm_in_cnsi_biwt;
  wire plm_in_cnsi_bdwt;
  wire plm_in_cnsi_we_d_load_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cnsi_1_plm_in_cns_wait_ctrl
      softmax_sysc_load_load_plm_in_cnsi_1_plm_in_cns_wait_ctrl_inst (
      .load_wen(load_wen),
      .load_wten(load_wten),
      .plm_in_cnsi_oswt_unreg(plm_in_cnsi_oswt_unreg),
      .plm_in_cnsi_iswt0(plm_in_cnsi_iswt0),
      .plm_in_cnsi_biwt(plm_in_cnsi_biwt),
      .plm_in_cnsi_bdwt(plm_in_cnsi_bdwt),
      .plm_in_cnsi_we_d_load_sct_pff(plm_in_cnsi_we_d_load_sct_iff),
      .plm_in_cnsi_iswt0_pff(plm_in_cnsi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cnsi_1_plm_in_cns_wait_dp softmax_sysc_load_load_plm_in_cnsi_1_plm_in_cns_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cnsi_bawt(plm_in_cnsi_bawt),
      .plm_in_cnsi_biwt(plm_in_cnsi_biwt),
      .plm_in_cnsi_bdwt(plm_in_cnsi_bdwt)
    );
  assign plm_in_cnsi_we_d_pff = plm_in_cnsi_we_d_load_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_input_ready_req_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_input_ready_req_mioi (
  clk, rst, input_ready_req_req, input_ready_ack_ack, load_wen, load_wten, input_ready_req_mioi_oswt_unreg,
      input_ready_req_mioi_bawt, input_ready_req_mioi_iswt0, input_ready_req_mioi_wen_comp,
      input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_psct, input_ready_req_mioi_iswt0_pff
);
  input clk;
  input rst;
  output input_ready_req_req;
  input input_ready_ack_ack;
  input load_wen;
  input load_wten;
  input input_ready_req_mioi_oswt_unreg;
  output input_ready_req_mioi_bawt;
  input input_ready_req_mioi_iswt0;
  output input_ready_req_mioi_wen_comp;
  input input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_psct;
  input input_ready_req_mioi_iswt0_pff;


  // Interconnect Declarations
  wire input_ready_req_mioi_biwt;
  wire input_ready_req_mioi_bdwt;
  wire input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_sct;
  wire input_ready_req_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_handshake_t_req  input_ready_req_mioi (
      .this_req_req(input_ready_req_req),
      .this_ack_ack(input_ready_ack_ack),
      .ccs_ccore_start_rsc_dat(input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_sct),
      .ccs_ccore_done_sync_vld(input_ready_req_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_input_ready_req_mioi_input_ready_req_mio_wait_ctrl
      softmax_sysc_load_load_input_ready_req_mioi_input_ready_req_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .load_wen(load_wen),
      .load_wten(load_wten),
      .input_ready_req_mioi_oswt_unreg(input_ready_req_mioi_oswt_unreg),
      .input_ready_req_mioi_iswt0(input_ready_req_mioi_iswt0),
      .input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_psct(input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_psct),
      .input_ready_req_mioi_biwt(input_ready_req_mioi_biwt),
      .input_ready_req_mioi_bdwt(input_ready_req_mioi_bdwt),
      .input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_sct(input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_sct),
      .input_ready_req_mioi_ccs_ccore_done_sync_vld(input_ready_req_mioi_ccs_ccore_done_sync_vld),
      .input_ready_req_mioi_iswt0_pff(input_ready_req_mioi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_input_ready_req_mioi_input_ready_req_mio_wait_dp
      softmax_sysc_load_load_input_ready_req_mioi_input_ready_req_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_ready_req_mioi_oswt_unreg(input_ready_req_mioi_oswt_unreg),
      .input_ready_req_mioi_bawt(input_ready_req_mioi_bawt),
      .input_ready_req_mioi_wen_comp(input_ready_req_mioi_wen_comp),
      .input_ready_req_mioi_biwt(input_ready_req_mioi_biwt),
      .input_ready_req_mioi_bdwt(input_ready_req_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_chnl_Pop_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_chnl_Pop_mioi (
  clk, rst, dma_read_chnl_val, dma_read_chnl_rdy, dma_read_chnl_msg, load_wen, load_wten,
      dma_read_chnl_Pop_mioi_oswt_unreg, dma_read_chnl_Pop_mioi_bawt, dma_read_chnl_Pop_mioi_iswt0,
      dma_read_chnl_Pop_mioi_wen_comp, dma_read_chnl_Pop_mioi_return_rsc_z_mxwt,
      dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_psct, dma_read_chnl_Pop_mioi_iswt0_pff
);
  input clk;
  input rst;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  input load_wen;
  input load_wten;
  input dma_read_chnl_Pop_mioi_oswt_unreg;
  output dma_read_chnl_Pop_mioi_bawt;
  input dma_read_chnl_Pop_mioi_iswt0;
  output dma_read_chnl_Pop_mioi_wen_comp;
  output [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt;
  input dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_psct;
  input dma_read_chnl_Pop_mioi_iswt0_pff;


  // Interconnect Declarations
  wire [63:0] dma_read_chnl_Pop_mioi_return_rsc_z;
  wire dma_read_chnl_Pop_mioi_biwt;
  wire dma_read_chnl_Pop_mioi_bdwt;
  wire dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_sct;
  wire dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld;
  wire [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_Connections_InBlocking_dma_data_t_Connections_SYN_PORT_Pop
      dma_read_chnl_Pop_mioi (
      .this_val(dma_read_chnl_val),
      .this_rdy(dma_read_chnl_rdy),
      .this_msg(dma_read_chnl_msg),
      .return_rsc_z(dma_read_chnl_Pop_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_sct),
      .ccs_ccore_done_sync_vld(dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl
      softmax_sysc_load_load_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .load_wen(load_wen),
      .load_wten(load_wten),
      .dma_read_chnl_Pop_mioi_oswt_unreg(dma_read_chnl_Pop_mioi_oswt_unreg),
      .dma_read_chnl_Pop_mioi_iswt0(dma_read_chnl_Pop_mioi_iswt0),
      .dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_psct(dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_psct),
      .dma_read_chnl_Pop_mioi_biwt(dma_read_chnl_Pop_mioi_biwt),
      .dma_read_chnl_Pop_mioi_bdwt(dma_read_chnl_Pop_mioi_bdwt),
      .dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_sct(dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_sct),
      .dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld(dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld),
      .dma_read_chnl_Pop_mioi_iswt0_pff(dma_read_chnl_Pop_mioi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp
      softmax_sysc_load_load_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_chnl_Pop_mioi_oswt_unreg(dma_read_chnl_Pop_mioi_oswt_unreg),
      .dma_read_chnl_Pop_mioi_bawt(dma_read_chnl_Pop_mioi_bawt),
      .dma_read_chnl_Pop_mioi_wen_comp(dma_read_chnl_Pop_mioi_wen_comp),
      .dma_read_chnl_Pop_mioi_return_rsc_z_mxwt(dma_read_chnl_Pop_mioi_return_rsc_z_mxwt_pconst),
      .dma_read_chnl_Pop_mioi_return_rsc_z(dma_read_chnl_Pop_mioi_return_rsc_z),
      .dma_read_chnl_Pop_mioi_biwt(dma_read_chnl_Pop_mioi_biwt),
      .dma_read_chnl_Pop_mioi_bdwt(dma_read_chnl_Pop_mioi_bdwt)
    );
  assign dma_read_chnl_Pop_mioi_return_rsc_z_mxwt = dma_read_chnl_Pop_mioi_return_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_ctrl_Push_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_ctrl_Push_mioi (
  clk, rst, dma_read_ctrl_val, dma_read_ctrl_rdy, dma_read_ctrl_msg, load_wen, dma_read_ctrl_Push_mioi_m_index_rsc_dat,
      dma_read_ctrl_Push_mioi_oswt_unreg, dma_read_ctrl_Push_mioi_bawt, dma_read_ctrl_Push_mioi_iswt0,
      load_wten, dma_read_ctrl_Push_mioi_wen_comp, dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_psct,
      dma_read_ctrl_Push_mioi_iswt0_pff
);
  input clk;
  input rst;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  input load_wen;
  input [31:0] dma_read_ctrl_Push_mioi_m_index_rsc_dat;
  input dma_read_ctrl_Push_mioi_oswt_unreg;
  output dma_read_ctrl_Push_mioi_bawt;
  input dma_read_ctrl_Push_mioi_iswt0;
  input load_wten;
  output dma_read_ctrl_Push_mioi_wen_comp;
  input dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_psct;
  input dma_read_ctrl_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire dma_read_ctrl_Push_mioi_biwt;
  wire dma_read_ctrl_Push_mioi_bdwt;
  wire dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_sct;
  wire dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_dma_read_ctrl_Push_mioi_m_index_rsc_dat;
  assign nl_dma_read_ctrl_Push_mioi_m_index_rsc_dat = {21'b000000000000000000000
      , (dma_read_ctrl_Push_mioi_m_index_rsc_dat[10:7]) , 7'b0000000};
  esp_acc_softmax_sysc_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push
      dma_read_ctrl_Push_mioi (
      .this_val(dma_read_ctrl_val),
      .this_rdy(dma_read_ctrl_rdy),
      .this_msg(dma_read_ctrl_msg),
      .m_index_rsc_dat(nl_dma_read_ctrl_Push_mioi_m_index_rsc_dat[31:0]),
      .ccs_ccore_start_rsc_dat(dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_sct),
      .ccs_ccore_done_sync_vld(dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl
      softmax_sysc_load_load_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .load_wen(load_wen),
      .dma_read_ctrl_Push_mioi_oswt_unreg(dma_read_ctrl_Push_mioi_oswt_unreg),
      .dma_read_ctrl_Push_mioi_iswt0(dma_read_ctrl_Push_mioi_iswt0),
      .load_wten(load_wten),
      .dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_psct(dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_psct),
      .dma_read_ctrl_Push_mioi_biwt(dma_read_ctrl_Push_mioi_biwt),
      .dma_read_ctrl_Push_mioi_bdwt(dma_read_ctrl_Push_mioi_bdwt),
      .dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_sct(dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_sct),
      .dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld(dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .dma_read_ctrl_Push_mioi_iswt0_pff(dma_read_ctrl_Push_mioi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp
      softmax_sysc_load_load_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_ctrl_Push_mioi_oswt_unreg(dma_read_ctrl_Push_mioi_oswt_unreg),
      .dma_read_ctrl_Push_mioi_bawt(dma_read_ctrl_Push_mioi_bawt),
      .dma_read_ctrl_Push_mioi_wen_comp(dma_read_ctrl_Push_mioi_wen_comp),
      .dma_read_ctrl_Push_mioi_biwt(dma_read_ctrl_Push_mioi_biwt),
      .dma_read_ctrl_Push_mioi_bdwt(dma_read_ctrl_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_config
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_config (
  clk, rst, conf_done, done
);
  input clk;
  input rst;
  input conf_done;
  output done;
  reg done;


  // Interconnect Declarations
  wire [2:0] fsm_output;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_softmax_sysc_config_config_fsm_inst_CONFIG_LOOP_C_0_tr0;
  assign nl_softmax_sysc_config_config_fsm_inst_CONFIG_LOOP_C_0_tr0 = ~ conf_done;
  esp_acc_softmax_sysc_softmax_sysc_config_config_fsm softmax_sysc_config_config_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .CONFIG_LOOP_C_0_tr0(nl_softmax_sysc_config_config_fsm_inst_CONFIG_LOOP_C_0_tr0[0:0])
    );
  always @(posedge clk) begin
    if ( ~ rst ) begin
      done <= 1'b0;
    end
    else if ( conf_done & (fsm_output[1]) ) begin
      done <= 1'b1;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store_store
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store_store (
  clk, rst, conf_info, acc_done, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg,
      dma_write_chnl_val, dma_write_chnl_rdy, dma_write_chnl_msg, done, output_ready_req_req,
      output_ready_ack_ack, plm_out_cns_req_vz, plm_out_cns_rls_lz, plm_out_cnsi_q_d,
      plm_out_cnsi_radr_d, plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d
);
  input clk;
  input rst;
  input [31:0] conf_info;
  output acc_done;
  reg acc_done;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;
  input done;
  input output_ready_req_req;
  output output_ready_ack_ack;
  input plm_out_cns_req_vz;
  output plm_out_cns_rls_lz;
  input [31:0] plm_out_cnsi_q_d;
  output [6:0] plm_out_cnsi_radr_d;
  output plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations
  wire store_wen;
  wire output_ready_ack_mioi_bawt;
  reg output_ready_ack_mioi_iswt0;
  wire store_wten;
  wire output_ready_ack_mioi_wen_comp;
  reg output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_psct;
  wire dma_write_ctrl_Push_mioi_bawt;
  wire dma_write_ctrl_Push_mioi_wen_comp;
  reg dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct;
  wire dma_write_chnl_Push_mioi_bawt;
  wire dma_write_chnl_Push_mioi_wen_comp;
  reg dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct;
  wire plm_out_cnsi_bawt;
  wire [31:0] plm_out_cnsi_q_d_mxwt;
  wire plm_out_cns_rls_obj_bawt;
  wire plm_out_cns_req_obj_bawt;
  reg plm_out_cns_req_obj_iswt0;
  wire plm_out_cns_req_obj_wen_comp;
  reg [24:0] dma_write_ctrl_Push_mioi_m_index_rsc_dat_31_7;
  reg [31:0] dma_write_chnl_Push_mioi_m_rsc_dat_31_0;
  wire [6:0] fsm_output;
  wire [4:0] STORE_BATCH_LOOP_acc_3_tmp;
  wire [5:0] nl_STORE_BATCH_LOOP_acc_3_tmp;
  wire [7:0] STORE_LOOP_acc_2_tmp;
  wire [8:0] nl_STORE_LOOP_acc_2_tmp;
  wire STORE_BATCH_LOOP_and_12_tmp;
  wire STORE_BATCH_LOOP_and_8_tmp;
  wire or_dcpl_6;
  wire and_dcpl_2;
  wire or_tmp_10;
  wire and_dcpl_12;
  wire or_dcpl_23;
  wire and_dcpl_14;
  wire and_dcpl_16;
  wire or_dcpl_25;
  wire or_dcpl_27;
  wire or_dcpl_28;
  wire and_dcpl_21;
  wire and_dcpl_23;
  wire and_dcpl_24;
  wire or_dcpl_34;
  wire and_dcpl_25;
  wire and_dcpl_34;
  wire and_dcpl_35;
  wire and_dcpl_40;
  wire or_tmp_48;
  wire mux_tmp_58;
  wire and_dcpl_42;
  wire or_dcpl_38;
  wire or_dcpl_46;
  wire or_tmp_52;
  wire mux_tmp_61;
  wire or_dcpl_62;
  wire and_dcpl_69;
  wire and_tmp_14;
  wire and_dcpl_82;
  wire or_tmp_61;
  wire or_tmp_62;
  wire or_tmp_65;
  wire or_tmp_68;
  reg exitL_exit_STORE_LOOP_sva;
  wire STORE_BATCH_LOOP_nand_12_cse_1;
  reg exit_STORE_BATCH_LOOP_sva_1_st_2;
  reg STORE_LOOP_asn_itm_2;
  reg STORE_BATCH_LOOP_stage_v_2;
  reg STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_3;
  reg STORE_BATCH_LOOP_stage_v_3;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_st_4;
  reg STORE_BATCH_LOOP_stage_v_4;
  reg exit_STORE_BATCH_LOOP_sva_1_st_1;
  reg STORE_LOOP_asn_itm_1;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_st_1;
  reg STORE_BATCH_LOOP_stage_0_3;
  reg STORE_BATCH_LOOP_stage_0_4;
  reg STORE_LOOP_asn_itm;
  reg STORE_BATCH_LOOP_stage_0;
  reg STORE_BATCH_LOOP_stage_0_2;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_st_2;
  reg STORE_BATCH_LOOP_stage_0_1;
  reg STORE_BATCH_LOOP_stage_v;
  reg STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_2;
  reg reg_output_ready_ack_mioi_oswt_cse;
  reg reg_dma_write_chnl_Push_mioi_iswt0_cse;
  reg reg_plm_out_cnsi_iswt0_cse;
  reg reg_plm_out_cns_rls_obj_iswt0_cse;
  wire and_230_cse;
  wire STORE_BATCH_LOOP_and_14_cse;
  wire nand_16_cse;
  wire or_18_cse;
  wire nor_cse;
  wire and_233_cse;
  wire ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_and_cse;
  reg [6:0] plm_out_cnsi_radr_d_reg;
  wire [6:0] STORE_LOOP_i_mux_rmff;
  wire plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_reg;
  wire and_127_rmff;
  wire and_121_rmff;
  wire softmax_sysc_store_compute_handshake_softmax_sysc_store_compute_handshake_or_rmff;
  wire [24:0] STORE_BATCH_LOOP_mux_rmff;
  wire STORE_BATCH_LOOP_STORE_BATCH_LOOP_or_5_rmff;
  wire [31:0] STORE_LOOP_data_mux_rmff;
  wire STORE_LOOP_STORE_LOOP_or_rmff;
  reg [31:0] config_batch_sva;
  reg STORE_BATCH_LOOP_stage_v_1;
  reg exit_STORE_BATCH_LOOP_sva_1_st;
  reg STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm;
  reg [24:0] STORE_BATCH_LOOP_acc_4_itm_1;
  reg [6:0] STORE_LOOP_i_slc_STORE_LOOP_i_7_0_6_0_itm_1;
  reg [6:0] STORE_LOOP_i_slc_STORE_LOOP_i_7_0_6_0_itm_2;
  reg STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_1;
  reg [6:0] STORE_LOOP_i_7_0_lpi_1_6_0;
  reg [3:0] STORE_BATCH_LOOP_b_4_0_sva_3_0;
  wire exitL_exit_STORE_LOOP_sva_mx1w0;
  wire STORE_BATCH_LOOP_stage_v_2_mx0c1;
  wire STORE_BATCH_LOOP_stage_0_3_mx0c1;
  wire STORE_BATCH_LOOP_or_1_cse_1;
  wire STORE_BATCH_LOOP_or_2_cse_1;
  wire STORE_BATCH_LOOP_STORE_BATCH_LOOP_or_cse_1;
  wire and_101_rgt;
  wire STORE_LOOP_i_and_6_itm;
  wire STORE_BATCH_LOOP_acc_1_itm_32_1;

  wire[0:0] or_142_nl;
  wire[0:0] or_146_nl;
  wire[0:0] or_150_nl;
  wire[3:0] STORE_BATCH_LOOP_b_mux_nl;
  wire[0:0] STORE_BATCH_LOOP_b_and_nl;
  wire[0:0] STORE_BATCH_LOOP_mux1h_nl;
  wire[0:0] and_78_nl;
  wire[0:0] and_80_nl;
  wire[0:0] or_111_nl;
  wire[0:0] STORE_BATCH_LOOP_mux_30_nl;
  wire[0:0] or_113_nl;
  wire[0:0] mux_70_nl;
  wire[0:0] or_118_nl;
  wire[0:0] or_124_nl;
  wire[24:0] STORE_BATCH_LOOP_acc_4_nl;
  wire[25:0] nl_STORE_BATCH_LOOP_acc_4_nl;
  wire[0:0] STORE_BATCH_LOOP_and_23_nl;
  wire[0:0] and_96_nl;
  wire[0:0] and_97_nl;
  wire[0:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_nl;
  wire[0:0] STORE_BATCH_LOOP_mux_29_nl;
  wire[0:0] nor_42_nl;
  wire[0:0] STORE_BATCH_LOOP_mux_28_nl;
  wire[0:0] or_120_nl;
  wire[0:0] mux_73_nl;
  wire[0:0] mux_72_nl;
  wire[0:0] mux_71_nl;
  wire[0:0] and_103_nl;
  wire[32:0] STORE_BATCH_LOOP_acc_1_nl;
  wire[33:0] nl_STORE_BATCH_LOOP_acc_1_nl;
  wire[6:0] STORE_LOOP_mux_6_nl;
  wire[0:0] and_57_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_softmax_sysc_store_store_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat;
  assign nl_softmax_sysc_store_store_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat
      = {STORE_BATCH_LOOP_mux_rmff , 7'b0000000};
  wire [63:0] nl_softmax_sysc_store_store_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_m_rsc_dat;
  assign nl_softmax_sysc_store_store_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_m_rsc_dat
      = {32'b11011110101011011011111011101111 , STORE_LOOP_data_mux_rmff};
  wire [0:0] nl_softmax_sysc_store_store_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_oswt_unreg;
  assign nl_softmax_sysc_store_store_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_oswt_unreg
      = and_dcpl_34 & (fsm_output[1]);
  wire [0:0] nl_softmax_sysc_store_store_plm_out_cns_rls_obj_inst_plm_out_cns_rls_obj_oswt_unreg;
  assign nl_softmax_sysc_store_store_plm_out_cns_rls_obj_inst_plm_out_cns_rls_obj_oswt_unreg
      = or_dcpl_25 & plm_out_cnsi_bawt & plm_out_cns_rls_obj_bawt & STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_3
      & (~ exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3) & and_dcpl_35 & (fsm_output[1]);
  wire [0:0] nl_softmax_sysc_store_store_store_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  assign nl_softmax_sysc_store_store_store_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0
      = ~ done;
  wire [0:0] nl_softmax_sysc_store_store_store_fsm_inst_STORE_BATCH_LOOP_C_0_tr0;
  assign nl_softmax_sysc_store_store_store_fsm_inst_STORE_BATCH_LOOP_C_0_tr0 = ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_and_cse
      | nor_cse | (~ STORE_BATCH_LOOP_stage_v_4) | STORE_BATCH_LOOP_stage_0_4 | STORE_BATCH_LOOP_stage_0_2
      | STORE_BATCH_LOOP_stage_0_1 | STORE_BATCH_LOOP_stage_0_3;
  esp_acc_softmax_sysc_softmax_sysc_store_store_output_ready_ack_mioi softmax_sysc_store_store_output_ready_ack_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .output_ready_req_req(output_ready_req_req),
      .output_ready_ack_ack(output_ready_ack_ack),
      .store_wen(store_wen),
      .output_ready_ack_mioi_oswt_unreg(or_tmp_61),
      .output_ready_ack_mioi_bawt(output_ready_ack_mioi_bawt),
      .output_ready_ack_mioi_iswt0(output_ready_ack_mioi_iswt0),
      .store_wten(store_wten),
      .output_ready_ack_mioi_wen_comp(output_ready_ack_mioi_wen_comp),
      .output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_psct(softmax_sysc_store_compute_handshake_softmax_sysc_store_compute_handshake_or_rmff),
      .output_ready_ack_mioi_iswt0_pff(or_tmp_65)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_ctrl_Push_mioi softmax_sysc_store_store_dma_write_ctrl_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_ctrl_val(dma_write_ctrl_val),
      .dma_write_ctrl_rdy(dma_write_ctrl_rdy),
      .dma_write_ctrl_msg(dma_write_ctrl_msg),
      .store_wen(store_wen),
      .store_wten(store_wten),
      .dma_write_ctrl_Push_mioi_m_index_rsc_dat(nl_softmax_sysc_store_store_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat[31:0]),
      .dma_write_ctrl_Push_mioi_oswt_unreg(and_121_rmff),
      .dma_write_ctrl_Push_mioi_bawt(dma_write_ctrl_Push_mioi_bawt),
      .dma_write_ctrl_Push_mioi_iswt0(reg_output_ready_ack_mioi_oswt_cse),
      .dma_write_ctrl_Push_mioi_wen_comp(dma_write_ctrl_Push_mioi_wen_comp),
      .dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct(STORE_BATCH_LOOP_STORE_BATCH_LOOP_or_5_rmff),
      .dma_write_ctrl_Push_mioi_iswt0_pff(or_tmp_61)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_dma_write_chnl_Push_mioi softmax_sysc_store_store_dma_write_chnl_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_chnl_val(dma_write_chnl_val),
      .dma_write_chnl_rdy(dma_write_chnl_rdy),
      .dma_write_chnl_msg(dma_write_chnl_msg),
      .store_wen(store_wen),
      .store_wten(store_wten),
      .dma_write_chnl_Push_mioi_m_rsc_dat(nl_softmax_sysc_store_store_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_m_rsc_dat[63:0]),
      .dma_write_chnl_Push_mioi_oswt_unreg(nl_softmax_sysc_store_store_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_oswt_unreg[0:0]),
      .dma_write_chnl_Push_mioi_bawt(dma_write_chnl_Push_mioi_bawt),
      .dma_write_chnl_Push_mioi_iswt0(reg_dma_write_chnl_Push_mioi_iswt0_cse),
      .dma_write_chnl_Push_mioi_wen_comp(dma_write_chnl_Push_mioi_wen_comp),
      .dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct(STORE_LOOP_STORE_LOOP_or_rmff),
      .dma_write_chnl_Push_mioi_iswt0_pff(or_tmp_68)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cnsi_1 softmax_sysc_store_store_plm_out_cnsi_1_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cnsi_q_d(plm_out_cnsi_q_d),
      .plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d(plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_reg),
      .store_wen(store_wen),
      .store_wten(store_wten),
      .plm_out_cnsi_oswt_unreg(or_tmp_68),
      .plm_out_cnsi_bawt(plm_out_cnsi_bawt),
      .plm_out_cnsi_iswt0(reg_plm_out_cnsi_iswt0_cse),
      .plm_out_cnsi_q_d_mxwt(plm_out_cnsi_q_d_mxwt),
      .plm_out_cnsi_iswt0_pff(and_127_rmff)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_rls_obj softmax_sysc_store_store_plm_out_cns_rls_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_rls_lz(plm_out_cns_rls_lz),
      .store_wen(store_wen),
      .store_wten(store_wten),
      .plm_out_cns_rls_obj_oswt_unreg(nl_softmax_sysc_store_store_plm_out_cns_rls_obj_inst_plm_out_cns_rls_obj_oswt_unreg[0:0]),
      .plm_out_cns_rls_obj_bawt(plm_out_cns_rls_obj_bawt),
      .plm_out_cns_rls_obj_iswt0(reg_plm_out_cns_rls_obj_iswt0_cse)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_plm_out_cns_req_obj softmax_sysc_store_store_plm_out_cns_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_req_vz(plm_out_cns_req_vz),
      .store_wen(store_wen),
      .plm_out_cns_req_obj_oswt_unreg(and_121_rmff),
      .plm_out_cns_req_obj_bawt(plm_out_cns_req_obj_bawt),
      .plm_out_cns_req_obj_iswt0(plm_out_cns_req_obj_iswt0),
      .plm_out_cns_req_obj_wen_comp(plm_out_cns_req_obj_wen_comp)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_staller softmax_sysc_store_store_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .store_wen(store_wen),
      .store_wten(store_wten),
      .output_ready_ack_mioi_wen_comp(output_ready_ack_mioi_wen_comp),
      .dma_write_ctrl_Push_mioi_wen_comp(dma_write_ctrl_Push_mioi_wen_comp),
      .dma_write_chnl_Push_mioi_wen_comp(dma_write_chnl_Push_mioi_wen_comp),
      .plm_out_cns_req_obj_wen_comp(plm_out_cns_req_obj_wen_comp)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store_store_fsm softmax_sysc_store_store_store_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .store_wen(store_wen),
      .fsm_output(fsm_output),
      .WAIT_FOR_CONFIG_LOOP_C_0_tr0(nl_softmax_sysc_store_store_store_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0[0:0]),
      .STORE_BATCH_LOOP_C_0_tr0(nl_softmax_sysc_store_store_store_fsm_inst_STORE_BATCH_LOOP_C_0_tr0[0:0])
    );
  assign and_121_rmff = and_dcpl_21 & and_dcpl_16 & and_dcpl_14 & STORE_BATCH_LOOP_stage_0_3
      & (fsm_output[1]);
  assign and_127_rmff = and_dcpl_42 & and_dcpl_40 & (~ exit_STORE_BATCH_LOOP_lpi_1_dfm_st_2)
      & (fsm_output[1]);
  assign or_142_nl = (~ (fsm_output[1])) | and_dcpl_23 | and_dcpl_24 | (~ plm_out_cnsi_bawt)
      | exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3 | or_dcpl_38;
  assign STORE_LOOP_data_mux_rmff = MUX_v_32_2_2(plm_out_cnsi_q_d_mxwt, dma_write_chnl_Push_mioi_m_rsc_dat_31_0,
      or_142_nl);
  assign STORE_LOOP_STORE_LOOP_or_rmff = (dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct
      & (~((or_dcpl_34 | exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3 | (~ STORE_BATCH_LOOP_stage_0_4)
      | (~ STORE_BATCH_LOOP_stage_v_3)) & and_dcpl_34 & (fsm_output[1])))) | or_tmp_68;
  assign or_146_nl = (~ (fsm_output[1])) | or_dcpl_23;
  assign STORE_BATCH_LOOP_mux_rmff = MUX_v_25_2_2(STORE_BATCH_LOOP_acc_4_itm_1, dma_write_ctrl_Push_mioi_m_index_rsc_dat_31_7,
      or_146_nl);
  assign STORE_BATCH_LOOP_STORE_BATCH_LOOP_or_5_rmff = (dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct
      & (~ or_tmp_62)) | or_tmp_61;
  assign or_150_nl = (~ (fsm_output[1])) | (~ mux_tmp_58) | and_dcpl_23 | or_dcpl_46
      | exit_STORE_BATCH_LOOP_lpi_1_dfm_st_2;
  assign STORE_LOOP_i_mux_rmff = MUX_v_7_2_2(STORE_LOOP_i_slc_STORE_LOOP_i_7_0_6_0_itm_2,
      plm_out_cnsi_radr_d_reg, or_150_nl);
  assign softmax_sysc_store_compute_handshake_softmax_sysc_store_compute_handshake_or_rmff
      = (output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_psct & (~(and_dcpl_12
      & (~(STORE_BATCH_LOOP_acc_1_itm_32_1 & STORE_LOOP_asn_itm & STORE_BATCH_LOOP_and_12_tmp))
      & (fsm_output[1])))) | or_tmp_65;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_and_cse
      = STORE_BATCH_LOOP_stage_0 & (and_dcpl_2 | (~ STORE_BATCH_LOOP_and_12_tmp));
  assign and_230_cse = (STORE_LOOP_acc_2_tmp[7]) & (STORE_BATCH_LOOP_acc_3_tmp[4]);
  assign STORE_BATCH_LOOP_and_14_cse = store_wen & (fsm_output[1]);
  assign or_18_cse = (~ STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_3) | plm_out_cns_rls_obj_bawt;
  assign and_233_cse = plm_out_cns_req_obj_bawt & dma_write_ctrl_Push_mioi_bawt;
  assign nand_16_cse = ~((STORE_BATCH_LOOP_acc_3_tmp[4]) & (STORE_LOOP_acc_2_tmp[7]));
  assign and_101_rgt = (~ exitL_exit_STORE_LOOP_sva) & STORE_BATCH_LOOP_and_12_tmp
      & (fsm_output[1]);
  assign STORE_LOOP_i_and_6_itm = STORE_BATCH_LOOP_and_14_cse & STORE_BATCH_LOOP_and_12_tmp;
  assign exitL_exit_STORE_LOOP_sva_mx1w0 = ~((STORE_BATCH_LOOP_acc_3_tmp[4]) | (~
      (STORE_LOOP_acc_2_tmp[7])));
  assign nl_STORE_BATCH_LOOP_acc_1_nl = ({29'b10000000000000000000000000000 , STORE_BATCH_LOOP_b_4_0_sva_3_0})
      + conv_u2u_32_33(~ config_batch_sva) + 33'b000000000000000000000000000000001;
  assign STORE_BATCH_LOOP_acc_1_nl = nl_STORE_BATCH_LOOP_acc_1_nl[32:0];
  assign STORE_BATCH_LOOP_acc_1_itm_32_1 = readslicef_33_1_32(STORE_BATCH_LOOP_acc_1_nl);
  assign nl_STORE_BATCH_LOOP_acc_3_tmp = conv_u2u_4_5(STORE_BATCH_LOOP_b_4_0_sva_3_0)
      + 5'b00001;
  assign STORE_BATCH_LOOP_acc_3_tmp = nl_STORE_BATCH_LOOP_acc_3_tmp[4:0];
  assign STORE_LOOP_mux_6_nl = MUX_v_7_2_2(STORE_LOOP_i_7_0_lpi_1_6_0, (signext_7_1(~
      STORE_BATCH_LOOP_acc_1_itm_32_1)), exitL_exit_STORE_LOOP_sva);
  assign nl_STORE_LOOP_acc_2_tmp = conv_u2u_7_8(STORE_LOOP_mux_6_nl) + 8'b00000001;
  assign STORE_LOOP_acc_2_tmp = nl_STORE_LOOP_acc_2_tmp[7:0];
  assign STORE_BATCH_LOOP_or_1_cse_1 = plm_out_cnsi_bawt | (~((~ exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3)
      & STORE_BATCH_LOOP_stage_v_3));
  assign STORE_BATCH_LOOP_or_2_cse_1 = plm_out_cns_rls_obj_bawt | (~(STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_3
      & (~ exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3) & STORE_BATCH_LOOP_stage_v_3));
  assign STORE_BATCH_LOOP_STORE_BATCH_LOOP_or_cse_1 = dma_write_chnl_Push_mioi_bawt
      | (~((~ exit_STORE_BATCH_LOOP_lpi_1_dfm_st_4) & STORE_BATCH_LOOP_stage_v_4));
  assign STORE_BATCH_LOOP_nand_12_cse_1 = ~((~ exit_STORE_BATCH_LOOP_sva_1_st_2)
      & STORE_LOOP_asn_itm_2 & STORE_BATCH_LOOP_stage_v_2);
  assign STORE_BATCH_LOOP_and_12_tmp = STORE_BATCH_LOOP_stage_v & (~(STORE_BATCH_LOOP_stage_v_1
      & (~ STORE_BATCH_LOOP_and_8_tmp))) & STORE_BATCH_LOOP_stage_0_1 & (dma_write_ctrl_Push_mioi_bawt
      | STORE_BATCH_LOOP_nand_12_cse_1) & (plm_out_cns_req_obj_bawt | STORE_BATCH_LOOP_nand_12_cse_1)
      & STORE_BATCH_LOOP_or_1_cse_1 & STORE_BATCH_LOOP_or_2_cse_1 & STORE_BATCH_LOOP_STORE_BATCH_LOOP_or_cse_1;
  assign STORE_BATCH_LOOP_and_8_tmp = STORE_BATCH_LOOP_stage_v_1 & (~(STORE_BATCH_LOOP_stage_v_2
      & or_dcpl_62)) & STORE_BATCH_LOOP_stage_0_2 & (output_ready_ack_mioi_bawt |
      (~((~ exit_STORE_BATCH_LOOP_sva_1_st_1) & STORE_LOOP_asn_itm_1))) & STORE_BATCH_LOOP_or_1_cse_1
      & STORE_BATCH_LOOP_or_2_cse_1 & STORE_BATCH_LOOP_STORE_BATCH_LOOP_or_cse_1;
  assign nor_cse = ~(exit_STORE_BATCH_LOOP_lpi_1_dfm_st_4 | dma_write_chnl_Push_mioi_bawt);
  assign or_dcpl_6 = STORE_BATCH_LOOP_acc_1_itm_32_1 | (~ exitL_exit_STORE_LOOP_sva);
  assign and_dcpl_2 = or_dcpl_6 & nand_16_cse;
  assign or_tmp_10 = exit_STORE_BATCH_LOOP_lpi_1_dfm_st_4 | dma_write_chnl_Push_mioi_bawt;
  assign and_dcpl_12 = (~ exit_STORE_BATCH_LOOP_sva_1_st_1) & STORE_LOOP_asn_itm_1
      & STORE_BATCH_LOOP_and_8_tmp;
  assign or_dcpl_23 = exit_STORE_BATCH_LOOP_sva_1_st_1 | (~ STORE_LOOP_asn_itm_1)
      | (~ STORE_BATCH_LOOP_and_8_tmp);
  assign and_dcpl_14 = STORE_LOOP_asn_itm_2 & STORE_BATCH_LOOP_stage_v_2;
  assign and_dcpl_16 = dma_write_ctrl_Push_mioi_bawt & plm_out_cns_req_obj_bawt &
      (~ exit_STORE_BATCH_LOOP_sva_1_st_2);
  assign or_dcpl_25 = or_tmp_10 | (~ STORE_BATCH_LOOP_stage_v_4);
  assign or_dcpl_27 = (or_18_cse & plm_out_cnsi_bawt) | exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3;
  assign or_dcpl_28 = ~((~(or_dcpl_27 & STORE_BATCH_LOOP_stage_0_4)) & STORE_BATCH_LOOP_stage_v_3);
  assign and_dcpl_21 = or_dcpl_28 & or_dcpl_25;
  assign and_dcpl_23 = nor_cse & STORE_BATCH_LOOP_stage_v_4;
  assign and_dcpl_24 = (~ plm_out_cns_rls_obj_bawt) & STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_3;
  assign or_dcpl_34 = and_dcpl_24 | (~ plm_out_cnsi_bawt);
  assign and_dcpl_25 = or_dcpl_34 & (~ exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3);
  assign and_dcpl_34 = (~ exit_STORE_BATCH_LOOP_lpi_1_dfm_st_4) & dma_write_chnl_Push_mioi_bawt
      & STORE_BATCH_LOOP_stage_v_4;
  assign and_dcpl_35 = STORE_BATCH_LOOP_stage_0_4 & STORE_BATCH_LOOP_stage_v_3;
  assign and_dcpl_40 = STORE_BATCH_LOOP_stage_v_2 & STORE_BATCH_LOOP_stage_0_3;
  assign or_tmp_48 = (~ STORE_LOOP_asn_itm_2) | exit_STORE_BATCH_LOOP_sva_1_st_2;
  assign and_57_nl = and_233_cse & or_dcpl_28;
  assign mux_tmp_58 = MUX_s_1_2_2(and_57_nl, or_dcpl_28, or_tmp_48);
  assign and_dcpl_42 = mux_tmp_58 & or_dcpl_25;
  assign or_dcpl_38 = ~(STORE_BATCH_LOOP_stage_0_4 & STORE_BATCH_LOOP_stage_v_3);
  assign or_dcpl_46 = ~(STORE_BATCH_LOOP_stage_v_2 & STORE_BATCH_LOOP_stage_0_3);
  assign or_tmp_52 = ~(nand_16_cse & or_dcpl_6);
  assign mux_tmp_61 = MUX_s_1_2_2(STORE_BATCH_LOOP_stage_v, or_tmp_52, STORE_BATCH_LOOP_and_12_tmp);
  assign or_dcpl_62 = (~ mux_tmp_58) | and_dcpl_23 | or_dcpl_46;
  assign and_dcpl_69 = and_dcpl_42 & and_dcpl_40;
  assign and_tmp_14 = and_dcpl_35 & or_dcpl_27;
  assign and_dcpl_82 = exitL_exit_STORE_LOOP_sva & STORE_BATCH_LOOP_and_12_tmp;
  assign or_tmp_61 = and_dcpl_12 & (fsm_output[1]);
  assign or_tmp_62 = and_dcpl_21 & and_dcpl_16 & and_dcpl_14 & or_dcpl_23 & STORE_BATCH_LOOP_stage_0_3
      & (fsm_output[1]);
  assign or_tmp_65 = STORE_BATCH_LOOP_acc_1_itm_32_1 & STORE_LOOP_asn_itm & STORE_BATCH_LOOP_and_12_tmp
      & (fsm_output[1]);
  assign or_tmp_68 = or_dcpl_25 & or_18_cse & plm_out_cnsi_bawt & (~ exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3)
      & and_dcpl_35 & (fsm_output[1]);
  assign STORE_BATCH_LOOP_stage_v_2_mx0c1 = STORE_BATCH_LOOP_and_8_tmp & (fsm_output[1]);
  assign STORE_BATCH_LOOP_stage_0_3_mx0c1 = (and_dcpl_69 | STORE_BATCH_LOOP_and_8_tmp)
      & (fsm_output[1]);
  assign plm_out_cnsi_radr_d = STORE_LOOP_i_mux_rmff;
  assign plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d = plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      acc_done <= 1'b0;
    end
    else if ( store_wen & ((fsm_output[2]) | (fsm_output[5])) ) begin
      acc_done <= ~ (fsm_output[5]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cns_req_obj_iswt0 <= 1'b0;
    end
    else if ( store_wen & (or_tmp_61 | or_tmp_62) ) begin
      plm_out_cns_req_obj_iswt0 <= ~ or_tmp_62;
    end
  end
  always @(posedge clk) begin
    if ( store_wen ) begin
      dma_write_chnl_Push_mioi_m_rsc_dat_31_0 <= STORE_LOOP_data_mux_rmff;
      dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct <= STORE_LOOP_STORE_LOOP_or_rmff;
      dma_write_ctrl_Push_mioi_m_index_rsc_dat_31_7 <= STORE_BATCH_LOOP_mux_rmff;
      dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_psct <= STORE_BATCH_LOOP_STORE_BATCH_LOOP_or_5_rmff;
      plm_out_cnsi_radr_d_reg <= STORE_LOOP_i_mux_rmff;
      output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_psct <= softmax_sysc_store_compute_handshake_softmax_sysc_store_compute_handshake_or_rmff;
      STORE_BATCH_LOOP_b_4_0_sva_3_0 <= MUX_v_4_2_2(4'b0000, STORE_BATCH_LOOP_b_mux_nl,
          (fsm_output[1]));
      config_batch_sva <= MUX_v_32_2_2(conf_info, config_batch_sva, fsm_output[1]);
      STORE_LOOP_i_slc_STORE_LOOP_i_7_0_6_0_itm_2 <= MUX_v_7_2_2(STORE_LOOP_i_slc_STORE_LOOP_i_7_0_6_0_itm_2,
          STORE_LOOP_i_slc_STORE_LOOP_i_7_0_6_0_itm_1, STORE_BATCH_LOOP_and_8_tmp);
      STORE_BATCH_LOOP_stage_v_1 <= ((STORE_BATCH_LOOP_stage_v_1 & (~ STORE_BATCH_LOOP_and_8_tmp))
          | STORE_BATCH_LOOP_and_12_tmp) & (fsm_output[1]);
      STORE_BATCH_LOOP_acc_4_itm_1 <= MUX_v_25_2_2(STORE_BATCH_LOOP_acc_4_itm_1,
          STORE_BATCH_LOOP_acc_4_nl, STORE_BATCH_LOOP_and_23_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_output_ready_ack_mioi_oswt_cse <= 1'b0;
      output_ready_ack_mioi_iswt0 <= 1'b0;
      reg_dma_write_chnl_Push_mioi_iswt0_cse <= 1'b0;
      reg_plm_out_cnsi_iswt0_cse <= 1'b0;
      reg_plm_out_cns_rls_obj_iswt0_cse <= 1'b0;
      STORE_BATCH_LOOP_stage_v <= 1'b0;
      STORE_BATCH_LOOP_stage_0 <= 1'b0;
      STORE_LOOP_asn_itm <= 1'b0;
      exitL_exit_STORE_LOOP_sva <= 1'b0;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_st_2 <= 1'b0;
      STORE_BATCH_LOOP_stage_v_3 <= 1'b0;
      STORE_BATCH_LOOP_stage_v_4 <= 1'b0;
      STORE_BATCH_LOOP_stage_0_1 <= 1'b0;
      STORE_BATCH_LOOP_stage_0_2 <= 1'b0;
      STORE_BATCH_LOOP_stage_0_4 <= 1'b0;
    end
    else if ( store_wen ) begin
      reg_output_ready_ack_mioi_oswt_cse <= or_tmp_61;
      output_ready_ack_mioi_iswt0 <= or_tmp_65;
      reg_dma_write_chnl_Push_mioi_iswt0_cse <= or_tmp_68;
      reg_plm_out_cnsi_iswt0_cse <= and_127_rmff;
      reg_plm_out_cns_rls_obj_iswt0_cse <= and_dcpl_42 & and_dcpl_40 & (~ exit_STORE_BATCH_LOOP_lpi_1_dfm_st_2)
          & STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_2 & (fsm_output[1]);
      STORE_BATCH_LOOP_stage_v <= ~((~(STORE_BATCH_LOOP_stage_v & (~(((~ or_dcpl_6)
          | and_230_cse | (~ STORE_BATCH_LOOP_stage_0)) & STORE_BATCH_LOOP_and_12_tmp))))
          & (~((~ mux_tmp_61) & STORE_BATCH_LOOP_stage_0)) & (fsm_output[1]));
      STORE_BATCH_LOOP_stage_0 <= ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_and_cse
          | (~ (fsm_output[1]));
      STORE_LOOP_asn_itm <= STORE_BATCH_LOOP_mux1h_nl | (~ (fsm_output[1]));
      exitL_exit_STORE_LOOP_sva <= STORE_BATCH_LOOP_mux_30_nl | (~ (fsm_output[1]));
      exit_STORE_BATCH_LOOP_lpi_1_dfm_st_2 <= MUX_s_1_2_2(exit_STORE_BATCH_LOOP_lpi_1_dfm_st_2,
          exit_STORE_BATCH_LOOP_lpi_1_dfm_st_1, STORE_BATCH_LOOP_and_8_tmp);
      STORE_BATCH_LOOP_stage_v_3 <= ((STORE_BATCH_LOOP_stage_v_3 & (~((~ mux_70_nl)
          & or_dcpl_25 & and_dcpl_35))) | and_dcpl_69) & (fsm_output[1]);
      STORE_BATCH_LOOP_stage_v_4 <= ((STORE_BATCH_LOOP_stage_v_4 & (~((and_dcpl_25
          | or_dcpl_38) & or_tmp_10))) | (or_dcpl_27 & or_dcpl_25 & and_dcpl_35))
          & (fsm_output[1]);
      STORE_BATCH_LOOP_stage_0_1 <= ~((~(ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_nl
          & (~(or_tmp_52 & STORE_BATCH_LOOP_and_12_tmp)))) & (fsm_output[1]));
      STORE_BATCH_LOOP_stage_0_2 <= STORE_BATCH_LOOP_mux_29_nl & (fsm_output[1]);
      STORE_BATCH_LOOP_stage_0_4 <= STORE_BATCH_LOOP_mux_28_nl & (fsm_output[1]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      STORE_BATCH_LOOP_stage_v_2 <= 1'b0;
    end
    else if ( store_wen & ((and_dcpl_42 & and_dcpl_40 & (~ STORE_BATCH_LOOP_and_8_tmp)
        & (fsm_output[1])) | (fsm_output[0]) | STORE_BATCH_LOOP_stage_v_2_mx0c1)
        ) begin
      STORE_BATCH_LOOP_stage_v_2 <= STORE_BATCH_LOOP_stage_v_2_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_STORE_BATCH_LOOP_sva_1_st_2 <= 1'b0;
      STORE_LOOP_asn_itm_2 <= 1'b0;
      STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_3 <= 1'b0;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3 <= 1'b0;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_st_4 <= 1'b0;
      exit_STORE_BATCH_LOOP_sva_1_st_1 <= 1'b0;
      STORE_LOOP_asn_itm_1 <= 1'b0;
    end
    else if ( STORE_BATCH_LOOP_and_14_cse ) begin
      exit_STORE_BATCH_LOOP_sva_1_st_2 <= MUX_s_1_2_2(exit_STORE_BATCH_LOOP_sva_1_st_2,
          exit_STORE_BATCH_LOOP_sva_1_st_1, STORE_BATCH_LOOP_and_8_tmp);
      STORE_LOOP_asn_itm_2 <= MUX_s_1_2_2(STORE_LOOP_asn_itm_2, STORE_LOOP_asn_itm_1,
          STORE_BATCH_LOOP_and_8_tmp);
      STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_3 <= MUX_s_1_2_2(STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_2,
          STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_3, or_dcpl_62);
      exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3 <= MUX_s_1_2_2(exit_STORE_BATCH_LOOP_lpi_1_dfm_st_2,
          exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3, or_dcpl_62);
      exit_STORE_BATCH_LOOP_lpi_1_dfm_st_4 <= MUX_s_1_2_2(exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3,
          exit_STORE_BATCH_LOOP_lpi_1_dfm_st_4, or_124_nl);
      exit_STORE_BATCH_LOOP_sva_1_st_1 <= MUX1HOT_s_1_3_2((~ STORE_BATCH_LOOP_acc_1_itm_32_1),
          exit_STORE_BATCH_LOOP_sva_1_st, exit_STORE_BATCH_LOOP_sva_1_st_1, {and_96_nl
          , and_97_nl , (~ STORE_BATCH_LOOP_and_12_tmp)});
      STORE_LOOP_asn_itm_1 <= MUX_s_1_2_2(STORE_LOOP_asn_itm_1, STORE_LOOP_asn_itm,
          STORE_BATCH_LOOP_and_12_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_2 <= 1'b0;
    end
    else if ( store_wen & STORE_BATCH_LOOP_and_8_tmp ) begin
      STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_2 <= STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( store_wen & (~((STORE_LOOP_acc_2_tmp[7]) | (~ STORE_BATCH_LOOP_and_12_tmp)))
        ) begin
      STORE_LOOP_i_7_0_lpi_1_6_0 <= STORE_LOOP_acc_2_tmp[6:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      STORE_BATCH_LOOP_stage_0_3 <= 1'b0;
    end
    else if ( store_wen & ((fsm_output[0]) | STORE_BATCH_LOOP_stage_0_3_mx0c1) )
        begin
      STORE_BATCH_LOOP_stage_0_3 <= STORE_BATCH_LOOP_stage_0_2 & STORE_BATCH_LOOP_stage_0_3_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_STORE_BATCH_LOOP_sva_1_st <= 1'b0;
    end
    else if ( store_wen & STORE_LOOP_asn_itm & STORE_BATCH_LOOP_and_12_tmp ) begin
      exit_STORE_BATCH_LOOP_sva_1_st <= ~ STORE_BATCH_LOOP_acc_1_itm_32_1;
    end
  end
  always @(posedge clk) begin
    if ( store_wen & ((and_dcpl_82 & (fsm_output[1])) | and_101_rgt) ) begin
      STORE_LOOP_i_slc_STORE_LOOP_i_7_0_6_0_itm_1 <= MUX_v_7_2_2((signext_7_1(~ STORE_BATCH_LOOP_acc_1_itm_32_1)),
          STORE_LOOP_i_7_0_lpi_1_6_0, and_101_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_1 <= 1'b0;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_st_1 <= 1'b0;
      STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm <= 1'b0;
    end
    else if ( STORE_LOOP_i_and_6_itm ) begin
      STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm_1 <= MUX_s_1_2_2((STORE_LOOP_acc_2_tmp[7]),
          STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm, and_103_nl);
      exit_STORE_BATCH_LOOP_lpi_1_dfm_st_1 <= (~ STORE_BATCH_LOOP_acc_1_itm_32_1)
          & exitL_exit_STORE_LOOP_sva;
      STORE_LOOP_i_slc_STORE_LOOP_i_7_0_7_itm <= STORE_LOOP_acc_2_tmp[7];
    end
  end
  assign STORE_BATCH_LOOP_b_and_nl = ((exitL_exit_STORE_LOOP_sva & (~ STORE_BATCH_LOOP_acc_1_itm_32_1)
      & STORE_LOOP_asn_itm) | (STORE_BATCH_LOOP_acc_3_tmp[4]) | (~ (STORE_LOOP_acc_2_tmp[7]))
      | (~ STORE_BATCH_LOOP_and_12_tmp)) & (fsm_output[1]);
  assign STORE_BATCH_LOOP_b_mux_nl = MUX_v_4_2_2((STORE_BATCH_LOOP_acc_3_tmp[3:0]),
      STORE_BATCH_LOOP_b_4_0_sva_3_0, STORE_BATCH_LOOP_b_and_nl);
  assign and_78_nl = and_dcpl_2 & STORE_BATCH_LOOP_stage_0 & STORE_BATCH_LOOP_and_12_tmp;
  assign and_80_nl = (~ STORE_BATCH_LOOP_stage_v) & STORE_BATCH_LOOP_stage_0;
  assign or_111_nl = mux_tmp_61 | (~ STORE_BATCH_LOOP_stage_0);
  assign STORE_BATCH_LOOP_mux1h_nl = MUX1HOT_s_1_3_2(exitL_exit_STORE_LOOP_sva_mx1w0,
      exitL_exit_STORE_LOOP_sva, STORE_LOOP_asn_itm, {and_78_nl , and_80_nl , or_111_nl});
  assign or_113_nl = (~ or_dcpl_6) | and_230_cse | (~ STORE_BATCH_LOOP_and_12_tmp);
  assign STORE_BATCH_LOOP_mux_30_nl = MUX_s_1_2_2(exitL_exit_STORE_LOOP_sva_mx1w0,
      exitL_exit_STORE_LOOP_sva, or_113_nl);
  assign or_118_nl = or_tmp_48 | and_233_cse | and_dcpl_25;
  assign mux_70_nl = MUX_s_1_2_2(and_dcpl_25, or_118_nl, and_dcpl_40);
  assign nl_STORE_BATCH_LOOP_acc_4_nl = (config_batch_sva[24:0]) + conv_u2u_4_25(STORE_BATCH_LOOP_b_4_0_sva_3_0);
  assign STORE_BATCH_LOOP_acc_4_nl = nl_STORE_BATCH_LOOP_acc_4_nl[24:0];
  assign STORE_BATCH_LOOP_and_23_nl = STORE_BATCH_LOOP_and_12_tmp & (fsm_output[1]);
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_nl
      = MUX_s_1_2_2(STORE_BATCH_LOOP_stage_0_1, STORE_BATCH_LOOP_stage_0, STORE_BATCH_LOOP_and_12_tmp);
  assign nor_42_nl = ~(STORE_BATCH_LOOP_and_8_tmp | STORE_BATCH_LOOP_and_12_tmp);
  assign STORE_BATCH_LOOP_mux_29_nl = MUX_s_1_2_2(STORE_BATCH_LOOP_stage_0_1, STORE_BATCH_LOOP_stage_0_2,
      nor_42_nl);
  assign mux_71_nl = MUX_s_1_2_2(and_tmp_14, or_dcpl_28, and_233_cse);
  assign mux_72_nl = MUX_s_1_2_2(mux_71_nl, or_dcpl_28, or_tmp_48);
  assign mux_73_nl = MUX_s_1_2_2(and_tmp_14, mux_72_nl, and_dcpl_40);
  assign or_120_nl = (~ mux_73_nl) | and_dcpl_23;
  assign STORE_BATCH_LOOP_mux_28_nl = MUX_s_1_2_2(STORE_BATCH_LOOP_stage_0_3, STORE_BATCH_LOOP_stage_0_4,
      or_120_nl);
  assign or_124_nl = and_dcpl_25 | and_dcpl_23 | or_dcpl_38;
  assign and_96_nl = STORE_LOOP_asn_itm & STORE_BATCH_LOOP_and_12_tmp;
  assign and_97_nl = (~ STORE_LOOP_asn_itm) & STORE_BATCH_LOOP_and_12_tmp;
  assign and_103_nl = (~ STORE_BATCH_LOOP_acc_1_itm_32_1) & and_dcpl_82;

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [24:0] MUX_v_25_2_2;
    input [24:0] input_0;
    input [24:0] input_1;
    input [0:0] sel;
    reg [24:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_25_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input [0:0] vector;
  begin
    signext_7_1= {{6{vector[0]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [24:0] conv_u2u_4_25 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_25 = {{21{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [32:0] conv_u2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_33 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute_compute
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute_compute (
  clk, rst, conf_info, done, input_ready_req_req, input_ready_ack_ack, output_ready_req_req,
      output_ready_ack_ack, plm_in_cns_req_vz, plm_in_cns_rls_lz, plm_out_cns_req_vz,
      plm_out_cns_rls_lz, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      plm_in_cnsi_q_d, plm_in_cnsi_radr_d, plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d,
      plm_out_cnsi_d_d, plm_out_cnsi_wadr_d, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff,
      plm_out_cnsi_we_d_pff
);
  input clk;
  input rst;
  input [31:0] conf_info;
  input done;
  input input_ready_req_req;
  output input_ready_ack_ack;
  output output_ready_req_req;
  input output_ready_ack_ack;
  input plm_in_cns_req_vz;
  output plm_in_cns_rls_lz;
  input plm_out_cns_req_vz;
  output plm_out_cns_rls_lz;
  output [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d;
  input [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d;
  output [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d;
  output [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] plm_in_cnsi_q_d;
  output [6:0] plm_in_cnsi_radr_d;
  output plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d;
  output [31:0] plm_out_cnsi_d_d;
  output [6:0] plm_out_cnsi_wadr_d;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff;
  output plm_out_cnsi_we_d_pff;


  // Interconnect Declarations
  wire compute_wen;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt;
  wire compute_wten;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt;
  wire input_ready_ack_mioi_bawt;
  reg input_ready_ack_mioi_iswt0;
  wire input_ready_ack_mioi_wen_comp;
  reg input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_psct;
  wire output_ready_req_mioi_bawt;
  wire output_ready_req_mioi_wen_comp;
  reg output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_psct;
  wire plm_in_cnsi_bawt;
  wire [31:0] plm_in_cnsi_q_d_mxwt;
  wire plm_out_cnsi_bawt;
  wire plm_out_cns_rls_obj_bawt;
  wire CALC_SOFTMAX_LOOP_mul_cmp_bawt;
  wire [31:0] CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt;
  wire plm_in_cns_rls_obj_bawt;
  wire plm_in_cns_req_obj_bawt;
  reg plm_in_cns_req_obj_iswt0;
  wire plm_in_cns_req_obj_wen_comp;
  wire plm_out_cns_req_obj_bawt;
  reg plm_out_cns_req_obj_iswt0;
  wire plm_out_cns_req_obj_wen_comp;
  wire [2:0] fsm_output;
  wire [7:0] CALC_SOFTMAX_LOOP_acc_1_tmp;
  wire [8:0] nl_CALC_SOFTMAX_LOOP_acc_1_tmp;
  wire COMPUTE_BATCH_LOOP_and_33_tmp;
  wire COMPUTE_BATCH_LOOP_and_28_tmp;
  wire COMPUTE_BATCH_LOOP_and_23_tmp;
  wire COMPUTE_BATCH_LOOP_and_19_tmp;
  wire [73:0] SUM_EXP_LOOP_acc_1_tmp;
  wire [74:0] nl_SUM_EXP_LOOP_acc_1_tmp;
  wire COMPUTE_BATCH_LOOP_and_16_tmp;
  wire COMPUTE_BATCH_LOOP_and_13_tmp;
  wire [7:0] SUM_EXP_LOOP_acc_2_tmp;
  wire [8:0] nl_SUM_EXP_LOOP_acc_2_tmp;
  wire [7:0] CALC_EXP_LOOP_acc_1_tmp;
  wire [8:0] nl_CALC_EXP_LOOP_acc_1_tmp;
  wire mux_tmp_1;
  wire or_tmp_20;
  wire mux_tmp_29;
  wire nor_tmp_12;
  wire and_dcpl_52;
  wire and_dcpl_54;
  wire mux_tmp_187;
  wire mux_tmp_190;
  wire and_dcpl_64;
  wire mux_tmp_191;
  wire or_tmp_152;
  wire and_dcpl_82;
  wire and_dcpl_84;
  wire and_dcpl_103;
  wire and_dcpl_106;
  wire and_tmp_54;
  wire or_dcpl_16;
  wire and_dcpl_121;
  wire nand_tmp_12;
  wire and_dcpl_125;
  wire or_dcpl_45;
  wire or_tmp_202;
  wire mux_tmp_229;
  wire mux_tmp_232;
  wire or_dcpl_50;
  wire and_dcpl_140;
  wire or_dcpl_52;
  wire and_dcpl_142;
  wire and_dcpl_144;
  wire and_tmp_85;
  wire or_dcpl_53;
  wire and_dcpl_147;
  wire or_dcpl_56;
  wire or_dcpl_57;
  wire and_dcpl_165;
  wire and_dcpl_166;
  wire and_dcpl_214;
  wire and_dcpl_220;
  wire and_dcpl_240;
  wire and_dcpl_243;
  wire and_dcpl_246;
  wire or_dcpl_140;
  wire and_dcpl_301;
  wire or_tmp_309;
  wire or_tmp_320;
  wire or_tmp_322;
  wire or_tmp_337;
  wire or_tmp_339;
  wire or_tmp_431;
  reg exitL_exit_CALC_SOFTMAX_LOOP_sva;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_st_8;
  reg CALC_SOFTMAX_LOOP_asn_itm_8;
  reg COMPUTE_BATCH_LOOP_stage_v_8;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_10;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_1;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1_mx1w0;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0_mx1w0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1;
  wire CALC_SOFTMAX_LOOP_and_4_ssc_1;
  wire CALC_SOFTMAX_LOOP_and_5_ssc_1;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0;
  wire CALC_SOFTMAX_LOOP_equal_tmp_2;
  wire CALC_EXP_LOOP_and_svs_1;
  wire CALC_SOFTMAX_LOOP_or_tmp_1;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_5;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_4;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1;
  reg COMPUTE_BATCH_LOOP_asn_2_itm_4;
  reg CALC_EXP_LOOP_and_svs_st_4;
  reg CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_4;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_2;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1;
  reg ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_itm_1;
  reg COMPUTE_BATCH_LOOP_asn_2_itm_5;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_3;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0;
  reg COMPUTE_BATCH_LOOP_stage_v_7;
  reg COMPUTE_BATCH_LOOP_stage_0_8;
  reg COMPUTE_BATCH_LOOP_stage_0_10;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0;
  reg COMPUTE_BATCH_LOOP_stage_0_9;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_7;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0;
  reg COMPUTE_BATCH_LOOP_stage_0;
  reg COMPUTE_BATCH_LOOP_stage_v;
  reg CALC_SOFTMAX_LOOP_asn_itm;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_0;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_10;
  reg COMPUTE_BATCH_LOOP_stage_0_6;
  reg CALC_SOFTMAX_LOOP_and_10_itm_5;
  reg CALC_SOFTMAX_LOOP_and_10_itm_4;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_0;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_1;
  reg CALC_SOFTMAX_LOOP_asn_itm_1;
  reg CALC_SOFTMAX_LOOP_asn_1_itm_1;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_2;
  reg CALC_SOFTMAX_LOOP_asn_itm_2;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_3;
  reg CALC_SOFTMAX_LOOP_asn_itm_3;
  reg CALC_SOFTMAX_LOOP_asn_1_itm_3;
  reg CALC_SOFTMAX_LOOP_asn_1_itm_2;
  reg COMPUTE_BATCH_LOOP_asn_2_itm_3;
  reg COMPUTE_BATCH_LOOP_stage_v_6;
  reg COMPUTE_BATCH_LOOP_stage_0_7;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_st_1;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_st_2;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_st_7;
  reg CALC_SOFTMAX_LOOP_asn_itm_7;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_8;
  reg CALC_EXP_LOOP_and_svs_st_3;
  reg CALC_EXP_LOOP_and_svs_st_2;
  reg reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_cse;
  reg reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_cse;
  reg reg_plm_in_cnsi_iswt0_cse;
  reg reg_plm_out_cnsi_iswt0_cse;
  reg reg_output_ready_req_mioi_iswt0_cse;
  reg reg_plm_out_cns_rls_obj_iswt0_cse;
  reg reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_1_cse;
  reg reg_plm_in_cns_rls_obj_iswt0_cse;
  wire CALC_SOFTMAX_LOOP_and_31_cse;
  wire COMPUTE_BATCH_LOOP_and_37_cse;
  wire and_826_cse;
  reg reg_COMPUTE_BATCH_LOOP_stage_v_3_cse;
  reg reg_COMPUTE_BATCH_LOOP_stage_v_5_cse;
  reg reg_COMPUTE_BATCH_LOOP_stage_v_9_cse;
  reg reg_COMPUTE_BATCH_LOOP_stage_v_10_cse;
  wire or_106_cse;
  wire or_cse;
  wire or_8_cse;
  wire or_107_cse;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_and_cse;
  wire nor_127_cse;
  wire or_181_cse;
  wire or_48_cse;
  wire or_46_cse;
  wire nor_129_cse;
  wire nor_3_cse;
  wire or_120_cse;
  wire mux_271_cse;
  wire nor_95_cse;
  wire mux_141_cse;
  wire and_23_cse;
  wire and_244_cse;
  wire mux_212_cse;
  wire mux_244_cse;
  wire mux_243_cse;
  wire mux_248_cse;
  wire mux_21_cse;
  wire and_226_cse;
  reg [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d_reg;
  wire [66:0] ac_math_ac_shift_left_21_1_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_1_rmff;
  reg [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d_reg;
  wire [6:0] CALC_SOFTMAX_LOOP_i_mux_1_rmff;
  reg [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d_reg;
  wire [6:0] CALC_EXP_LOOP_i_mux_rmff;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff;
  wire and_443_rmff;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  wire and_447_rmff;
  reg [6:0] plm_in_cnsi_radr_d_reg;
  wire [6:0] CALC_EXP_LOOP_i_mux_1_rmff;
  wire plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_reg;
  wire and_459_rmff;
  reg [31:0] plm_out_cnsi_d_d_reg;
  wire [31:0] CALC_SOFTMAX_LOOP_mux_1_rmff;
  reg [6:0] plm_out_cnsi_wadr_d_reg;
  wire [6:0] CALC_SOFTMAX_LOOP_i_mux_rmff;
  wire plm_out_cnsi_we_d_iff;
  wire and_463_rmff;
  wire and_445_rmff;
  wire softmax_sysc_compute_load_handshake_softmax_sysc_compute_load_handshake_or_rmff;
  wire softmax_sysc_compute_store_handshake_softmax_sysc_compute_store_handshake_or_rmff;
  reg [93:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1;
  reg [73:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_1_1;
  wire [73:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_mx1;
  wire and_837_tmp;
  wire [93:0] operator_94_21_false_AC_TRN_AC_WRAP_rshift_itm;
  wire [72:0] operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm;
  wire mux_291_itm;
  reg [73:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1;
  reg [31:0] config_batch_sva;
  reg [31:0] COMPUTE_BATCH_LOOP_b_sva;
  reg COMPUTE_BATCH_LOOP_stage_v_1;
  reg COMPUTE_BATCH_LOOP_stage_v_2;
  reg COMPUTE_BATCH_LOOP_stage_v_4;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_st;
  reg CALC_EXP_LOOP_and_svs_st;
  reg [10:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm;
  reg [9:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_9_0_itm;
  reg [7:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm;
  reg CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm;
  reg CALC_SOFTMAX_LOOP_and_10_itm;
  reg [10:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_itm_1;
  reg [9:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18_0_1_itm_1;
  reg [6:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_32_14_18_12_itm_1;
  reg [6:0] CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_1;
  reg [6:0] CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_2;
  reg [10:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm_1;
  reg [9:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_9_0_itm_1;
  reg [7:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm_1;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_1;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_2;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_3;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_4;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_1;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_2;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_3;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_4;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_5;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_6;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_7;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_8;
  reg CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_1;
  reg CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_2;
  reg CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_3;
  reg CALC_SOFTMAX_LOOP_and_10_itm_1;
  reg CALC_SOFTMAX_LOOP_and_10_itm_2;
  reg CALC_SOFTMAX_LOOP_and_10_itm_3;
  reg CALC_SOFTMAX_LOOP_asn_itm_4;
  reg CALC_SOFTMAX_LOOP_asn_itm_5;
  reg CALC_SOFTMAX_LOOP_asn_itm_6;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_st_3;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_st_4;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_st_5;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_st_6;
  reg CALC_EXP_LOOP_and_svs_st_1;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_6;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_1;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_2;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_3;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_4;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_5;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_6;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_7;
  reg COMPUTE_BATCH_LOOP_asn_2_itm_2;
  reg COMPUTE_BATCH_LOOP_stage_0_1;
  reg COMPUTE_BATCH_LOOP_stage_0_2;
  reg COMPUTE_BATCH_LOOP_stage_0_3;
  reg COMPUTE_BATCH_LOOP_stage_0_4;
  reg COMPUTE_BATCH_LOOP_stage_0_5;
  reg [6:0] CALC_EXP_LOOP_i_7_0_lpi_1_6_0;
  reg [6:0] SUM_EXP_LOOP_i_7_0_lpi_1_6_0;
  reg [6:0] CALC_SOFTMAX_LOOP_i_7_0_lpi_1_6_0;
  reg [6:0] CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_1_6_0;
  reg [6:0] CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_2_6_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0;
  wire plm_in_cns_req_obj_iswt0_mx0c1;
  wire plm_out_cns_req_obj_iswt0_mx0c1;
  wire COMPUTE_BATCH_LOOP_stage_0_mx1;
  wire exitL_exit_CALC_SOFTMAX_LOOP_sva_mx1w0;
  wire COMPUTE_BATCH_LOOP_stage_v_6_mx0c1;
  wire COMPUTE_BATCH_LOOP_stage_v_7_mx0c1;
  wire COMPUTE_BATCH_LOOP_stage_0_7_mx0c1;
  wire COMPUTE_BATCH_LOOP_stage_0_8_mx0c1;
  wire [10:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm_mx0w1;
  wire [11:0] nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm_mx0w1;
  wire [7:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm_mx0w1;
  wire [8:0] nl_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm_mx0w1;
  wire [66:0] operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1;
  wire COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_11_cse_1;
  wire COMPUTE_BATCH_LOOP_or_40_cse_1;
  wire COMPUTE_BATCH_LOOP_or_41_cse_1;
  wire COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_7_cse_1;
  wire COMPUTE_BATCH_LOOP_or_4_cse_1;
  wire COMPUTE_BATCH_LOOP_or_10_cse_1;
  wire COMPUTE_BATCH_LOOP_or_6_cse_1;
  wire COMPUTE_BATCH_LOOP_or_7_cse_1;
  wire COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_1_cse_1;
  wire CALC_SOFTMAX_LOOP_or_16_cse_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire [18:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire signed [19:0] nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire [6:0] libraries_leading_sign_74_0_cfd8a2a1b60025d53198d215150438e7bf24_1;
  wire CALC_EXP_LOOP_i_and_2_rgt;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_nand_1_cse;
  wire CALC_EXP_LOOP_i_and_4_cse;
  wire CALC_EXP_LOOP_i_and_3_cse;
  wire CALC_SOFTMAX_LOOP_and_72_cse;
  wire CALC_SOFTMAX_LOOP_and_74_cse;
  wire CALC_EXP_LOOP_and_6_cse;
  wire COMPUTE_BATCH_LOOP_and_64_cse;
  wire ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_and_cse;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_and_cse;
  wire CALC_EXP_LOOP_and_5_cse;
  wire CALC_SOFTMAX_LOOP_and_75_cse;
  wire COMPUTE_BATCH_LOOP_and_62_cse;
  wire CALC_SOFTMAX_LOOP_and_89_cse;
  wire COMPUTE_BATCH_LOOP_and_72_cse;
  wire CALC_SOFTMAX_LOOP_i_and_34_cse;
  wire CALC_SOFTMAX_LOOP_i_and_36_cse;
  wire COMPUTE_BATCH_LOOP_and_65_cse;
  wire CALC_SOFTMAX_LOOP_i_and_22_itm;
  wire CALC_EXP_LOOP_and_7_itm;
  wire COMPUTE_BATCH_LOOP_acc_itm_32_1;
  wire [18:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28;

  wire[0:0] or_482_nl;
  wire[0:0] or_483_nl;
  wire[0:0] mux_238_nl;
  wire[31:0] COMPUTE_BATCH_LOOP_b_mux_nl;
  wire[31:0] COMPUTE_BATCH_LOOP_acc_1_nl;
  wire[32:0] nl_COMPUTE_BATCH_LOOP_acc_1_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_b_and_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_mux1h_nl;
  wire[0:0] and_201_nl;
  wire[0:0] and_203_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_mux_86_nl;
  wire[0:0] or_240_nl;
  wire[0:0] and_228_nl;
  wire[0:0] and_227_nl;
  wire[0:0] mux_277_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] and_232_nl;
  wire[0:0] and_231_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] mux_293_nl;
  wire[0:0] mux_292_nl;
  wire[0:0] and_nl;
  wire[0:0] mux_302_nl;
  wire[0:0] and_810_nl;
  wire[10:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[2:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_2_nl;
  wire[6:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_3_nl;
  wire[0:0] and_284_nl;
  wire[0:0] and_285_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_i_and_17_nl;
  wire[0:0] operator_74_54_false_AC_TRN_AC_WRAP_1_mux_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_mux_85_nl;
  wire[0:0] nor_125_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_mux_84_nl;
  wire[0:0] nor_126_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_mux_83_nl;
  wire[0:0] nor_122_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_mux_82_nl;
  wire[0:0] nor_123_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_mux_81_nl;
  wire[0:0] nor_124_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] and_240_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_mux_80_nl;
  wire[0:0] mux_282_nl;
  wire[0:0] nor_94_nl;
  wire[0:0] mux_281_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_mux_79_nl;
  wire[0:0] mux_296_nl;
  wire[0:0] nand_20_nl;
  wire[0:0] mux_295_nl;
  wire[0:0] and_264_nl;
  wire[0:0] and_263_nl;
  wire[0:0] nand_21_nl;
  wire[0:0] and_375_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_24_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_2_nl;
  wire[9:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl;
  wire[0:0] and_371_nl;
  wire[0:0] and_372_nl;
  wire[0:0] or_444_nl;
  wire[32:0] COMPUTE_BATCH_LOOP_acc_nl;
  wire[33:0] nl_COMPUTE_BATCH_LOOP_acc_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_and_28_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_and_29_nl;
  wire[46:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl;
  wire signed [47:0] nl_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_7_nl;
  wire[2:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_1_nl;
  wire[6:0] CALC_SOFTMAX_LOOP_mux_112_nl;
  wire[6:0] CALC_SOFTMAX_LOOP_mux_111_nl;
  wire[7:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_3_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] or_634_nl;
  wire[0:0] mux_258_nl;
  wire[0:0] mux_256_nl;
  wire[0:0] nand_23_nl;
  wire[0:0] nor_1_nl;
  wire[0:0] and_111_nl;
  wire[0:0] and_110_nl;
  wire[0:0] mux_206_nl;
  wire[0:0] and_119_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] nor_98_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] mux_245_nl;
  wire[0:0] and_210_nl;
  wire[0:0] and_256_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] nor_78_nl;
  wire[0:0] or_154_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] nor_106_nl;
  wire[0:0] mux_269_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] and_225_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] and_813_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [73:0] nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_a;
  assign nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_a = {ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm_1
      , ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_9_0_itm_1
      , 53'b00000000000000000000000000000000000000000000000000000};
  wire [20:0] nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a = {ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_itm_1
      , ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18_0_1_itm_1};
  wire [72:0] nl_operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg_a = SUM_EXP_LOOP_acc_1_tmp[72:0];
  wire [0:0] nl_softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_inst_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg;
  assign nl_softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_inst_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg
      = (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_5) & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1)
      & COMPUTE_BATCH_LOOP_and_13_tmp & (fsm_output[1]);
  wire [0:0] nl_softmax_sysc_compute_compute_output_ready_req_mioi_inst_output_ready_req_mioi_oswt_unreg;
  assign nl_softmax_sysc_compute_compute_output_ready_req_mioi_inst_output_ready_req_mioi_oswt_unreg
      = and_dcpl_82 & (fsm_output[1]);
  wire [0:0] nl_softmax_sysc_compute_compute_plm_in_cnsi_1_inst_plm_in_cnsi_oswt_unreg;
  assign nl_softmax_sysc_compute_compute_plm_in_cnsi_1_inst_plm_in_cnsi_oswt_unreg
      = nor_127_cse & COMPUTE_BATCH_LOOP_and_19_tmp & (fsm_output[1]);
  wire [0:0] nl_softmax_sysc_compute_compute_plm_out_cnsi_1_inst_plm_out_cnsi_oswt_unreg;
  assign nl_softmax_sysc_compute_compute_plm_out_cnsi_1_inst_plm_out_cnsi_oswt_unreg
      = or_106_cse & or_181_cse & plm_out_cnsi_bawt & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0) & and_dcpl_84 & (fsm_output[1]);
  wire [93:0] nl_softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp_inst_CALC_SOFTMAX_LOOP_mul_cmp_b_compute;
  assign nl_softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp_inst_CALC_SOFTMAX_LOOP_mul_cmp_b_compute
      = ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1;
  wire [0:0] nl_softmax_sysc_compute_compute_plm_in_cns_rls_obj_inst_plm_in_cns_rls_obj_oswt_unreg;
  assign nl_softmax_sysc_compute_compute_plm_in_cns_rls_obj_inst_plm_in_cns_rls_obj_oswt_unreg
      = nor_127_cse & COMPUTE_BATCH_LOOP_and_19_tmp & CALC_EXP_LOOP_and_svs_st_3
      & (fsm_output[1]);
  wire [0:0] nl_softmax_sysc_compute_compute_plm_in_cns_req_obj_inst_plm_in_cns_req_obj_oswt_unreg;
  assign nl_softmax_sysc_compute_compute_plm_in_cns_req_obj_inst_plm_in_cns_req_obj_oswt_unreg
      = and_dcpl_54 & (fsm_output[1]);
  wire [0:0] nl_softmax_sysc_compute_compute_plm_out_cns_req_obj_inst_plm_out_cns_req_obj_oswt_unreg;
  assign nl_softmax_sysc_compute_compute_plm_out_cns_req_obj_inst_plm_out_cns_req_obj_oswt_unreg
      = and_tmp_54 & and_dcpl_64 & (fsm_output[1]);
  wire [0:0] nl_softmax_sysc_compute_compute_compute_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  assign nl_softmax_sysc_compute_compute_compute_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0
      = ~ done;
  wire [0:0] nl_softmax_sysc_compute_compute_compute_fsm_inst_COMPUTE_BATCH_LOOP_C_0_tr0;
  assign nl_softmax_sysc_compute_compute_compute_fsm_inst_COMPUTE_BATCH_LOOP_C_0_tr0
      = (~(reg_COMPUTE_BATCH_LOOP_stage_v_10_cse & (output_ready_req_mioi_bawt |
      (~(CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_10 & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_1
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_0) & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_10))))))
      | COMPUTE_BATCH_LOOP_stage_0_mx1 | COMPUTE_BATCH_LOOP_stage_0_1 | COMPUTE_BATCH_LOOP_stage_0_2
      | COMPUTE_BATCH_LOOP_stage_0_3 | COMPUTE_BATCH_LOOP_stage_0_4 | COMPUTE_BATCH_LOOP_stage_0_5
      | COMPUTE_BATCH_LOOP_stage_0_6 | COMPUTE_BATCH_LOOP_stage_0_7 | COMPUTE_BATCH_LOOP_stage_0_8
      | COMPUTE_BATCH_LOOP_stage_0_9 | COMPUTE_BATCH_LOOP_stage_0_10;
  esp_acc_softmax_sysc_mgc_shift_br_v5 #(.width_a(32'sd74),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd94)) operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_a[73:0]),
      .s(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm_1),
      .z(operator_94_21_false_AC_TRN_AC_WRAP_rshift_itm)
    );
  esp_acc_softmax_sysc_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd67)) operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_32_14_18_12_itm_1),
      .z(operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1)
    );
  esp_acc_softmax_sysc_mgc_shift_l_v5 #(.width_a(32'sd73),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd73)) operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg_a[72:0]),
      .s(libraries_leading_sign_74_0_cfd8a2a1b60025d53198d215150438e7bf24_1),
      .z(operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  esp_acc_softmax_sysc_leading_sign_74_0  leading_sign_74_0_rg (
      .mantissa(SUM_EXP_LOOP_acc_1_tmp),
      .rtn(libraries_leading_sign_74_0_cfd8a2a1b60025d53198d215150438e7bf24_1)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1
      softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg),
      .compute_wen(compute_wen),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg(nl_softmax_sysc_compute_compute_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_inst_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg[0:0]),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0(reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_cse),
      .compute_wten(compute_wten),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1(and_445_rmff),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1(reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_cse),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff(and_443_rmff),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff(and_447_rmff)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_input_ready_ack_mioi softmax_sysc_compute_compute_input_ready_ack_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .input_ready_req_req(input_ready_req_req),
      .input_ready_ack_ack(input_ready_ack_ack),
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .input_ready_ack_mioi_oswt_unreg(or_tmp_309),
      .input_ready_ack_mioi_bawt(input_ready_ack_mioi_bawt),
      .input_ready_ack_mioi_iswt0(input_ready_ack_mioi_iswt0),
      .input_ready_ack_mioi_wen_comp(input_ready_ack_mioi_wen_comp),
      .input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_psct(softmax_sysc_compute_load_handshake_softmax_sysc_compute_load_handshake_or_rmff),
      .input_ready_ack_mioi_iswt0_pff(or_tmp_320)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_output_ready_req_mioi softmax_sysc_compute_compute_output_ready_req_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .output_ready_req_req(output_ready_req_req),
      .output_ready_ack_ack(output_ready_ack_ack),
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .output_ready_req_mioi_oswt_unreg(nl_softmax_sysc_compute_compute_output_ready_req_mioi_inst_output_ready_req_mioi_oswt_unreg[0:0]),
      .output_ready_req_mioi_bawt(output_ready_req_mioi_bawt),
      .output_ready_req_mioi_iswt0(reg_output_ready_req_mioi_iswt0_cse),
      .output_ready_req_mioi_wen_comp(output_ready_req_mioi_wen_comp),
      .output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_psct(softmax_sysc_compute_store_handshake_softmax_sysc_compute_store_handshake_or_rmff),
      .output_ready_req_mioi_iswt0_pff(or_tmp_322)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cnsi_1 softmax_sysc_compute_compute_plm_in_cnsi_1_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cnsi_q_d(plm_in_cnsi_q_d),
      .plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d(plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_reg),
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .plm_in_cnsi_oswt_unreg(nl_softmax_sysc_compute_compute_plm_in_cnsi_1_inst_plm_in_cnsi_oswt_unreg[0:0]),
      .plm_in_cnsi_bawt(plm_in_cnsi_bawt),
      .plm_in_cnsi_iswt0(reg_plm_in_cnsi_iswt0_cse),
      .plm_in_cnsi_q_d_mxwt(plm_in_cnsi_q_d_mxwt),
      .plm_in_cnsi_iswt0_pff(and_459_rmff)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cnsi_1 softmax_sysc_compute_compute_plm_out_cnsi_1_inst
      (
      .clk(clk),
      .rst(rst),
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .plm_out_cnsi_oswt_unreg(nl_softmax_sysc_compute_compute_plm_out_cnsi_1_inst_plm_out_cnsi_oswt_unreg[0:0]),
      .plm_out_cnsi_bawt(plm_out_cnsi_bawt),
      .plm_out_cnsi_iswt0(reg_plm_out_cnsi_iswt0_cse),
      .plm_out_cnsi_we_d_pff(plm_out_cnsi_we_d_iff),
      .plm_out_cnsi_iswt0_pff(and_463_rmff)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_rls_obj softmax_sysc_compute_compute_plm_out_cns_rls_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_rls_lz(plm_out_cns_rls_lz),
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .plm_out_cns_rls_obj_oswt_unreg(or_tmp_322),
      .plm_out_cns_rls_obj_bawt(plm_out_cns_rls_obj_bawt),
      .plm_out_cns_rls_obj_iswt0(reg_plm_out_cns_rls_obj_iswt0_cse)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp_inst
      (
      .clk(clk),
      .rst(rst),
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg(and_463_rmff),
      .CALC_SOFTMAX_LOOP_mul_cmp_bawt(CALC_SOFTMAX_LOOP_mul_cmp_bawt),
      .CALC_SOFTMAX_LOOP_mul_cmp_iswt2(reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_1_cse),
      .CALC_SOFTMAX_LOOP_mul_cmp_a_compute(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt),
      .CALC_SOFTMAX_LOOP_mul_cmp_b_compute(nl_softmax_sysc_compute_compute_CALC_SOFTMAX_LOOP_mul_cmp_inst_CALC_SOFTMAX_LOOP_mul_cmp_b_compute[93:0]),
      .CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt(CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_rls_obj softmax_sysc_compute_compute_plm_in_cns_rls_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_rls_lz(plm_in_cns_rls_lz),
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .plm_in_cns_rls_obj_oswt_unreg(nl_softmax_sysc_compute_compute_plm_in_cns_rls_obj_inst_plm_in_cns_rls_obj_oswt_unreg[0:0]),
      .plm_in_cns_rls_obj_bawt(plm_in_cns_rls_obj_bawt),
      .plm_in_cns_rls_obj_iswt0(reg_plm_in_cns_rls_obj_iswt0_cse)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_in_cns_req_obj softmax_sysc_compute_compute_plm_in_cns_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_req_vz(plm_in_cns_req_vz),
      .compute_wen(compute_wen),
      .plm_in_cns_req_obj_oswt_unreg(nl_softmax_sysc_compute_compute_plm_in_cns_req_obj_inst_plm_in_cns_req_obj_oswt_unreg[0:0]),
      .plm_in_cns_req_obj_bawt(plm_in_cns_req_obj_bawt),
      .plm_in_cns_req_obj_iswt0(plm_in_cns_req_obj_iswt0),
      .plm_in_cns_req_obj_wen_comp(plm_in_cns_req_obj_wen_comp)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_plm_out_cns_req_obj softmax_sysc_compute_compute_plm_out_cns_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_req_vz(plm_out_cns_req_vz),
      .compute_wen(compute_wen),
      .plm_out_cns_req_obj_oswt_unreg(nl_softmax_sysc_compute_compute_plm_out_cns_req_obj_inst_plm_out_cns_req_obj_oswt_unreg[0:0]),
      .plm_out_cns_req_obj_bawt(plm_out_cns_req_obj_bawt),
      .plm_out_cns_req_obj_iswt0(plm_out_cns_req_obj_iswt0),
      .plm_out_cns_req_obj_wen_comp(plm_out_cns_req_obj_wen_comp)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_staller softmax_sysc_compute_compute_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .compute_wen(compute_wen),
      .compute_wten(compute_wten),
      .input_ready_ack_mioi_wen_comp(input_ready_ack_mioi_wen_comp),
      .output_ready_req_mioi_wen_comp(output_ready_req_mioi_wen_comp),
      .plm_in_cns_req_obj_wen_comp(plm_in_cns_req_obj_wen_comp),
      .plm_out_cns_req_obj_wen_comp(plm_out_cns_req_obj_wen_comp)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute_compute_fsm softmax_sysc_compute_compute_compute_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .compute_wen(compute_wen),
      .fsm_output(fsm_output),
      .WAIT_FOR_CONFIG_LOOP_C_0_tr0(nl_softmax_sysc_compute_compute_compute_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0[0:0]),
      .COMPUTE_BATCH_LOOP_C_0_tr0(nl_softmax_sysc_compute_compute_compute_fsm_inst_COMPUTE_BATCH_LOOP_C_0_tr0[0:0])
    );
  assign and_443_rmff = (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1) & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_4)
      & COMPUTE_BATCH_LOOP_and_16_tmp & (fsm_output[1]);
  assign and_445_rmff = (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_5) & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_0) & COMPUTE_BATCH_LOOP_and_13_tmp
      & (fsm_output[1]);
  assign and_447_rmff = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1 & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_4)
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0) & COMPUTE_BATCH_LOOP_and_16_tmp
      & (fsm_output[1]);
  assign and_459_rmff = nor_129_cse & COMPUTE_BATCH_LOOP_and_23_tmp & (fsm_output[1]);
  assign or_181_cse = plm_out_cns_rls_obj_bawt | (~ CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9);
  assign and_463_rmff = and_dcpl_106 & and_dcpl_103 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0)
      & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1 & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8)
      & COMPUTE_BATCH_LOOP_stage_v_8 & (fsm_output[1]);
  assign softmax_sysc_compute_store_handshake_softmax_sysc_compute_store_handshake_or_rmff
      = (output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_psct & (~(((~(plm_out_cnsi_bawt
      & plm_out_cns_rls_obj_bawt)) | (~(CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9
      & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1)) | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0
      | exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9 | or_dcpl_16) & and_dcpl_82 & (fsm_output[1]))))
      | or_tmp_322;
  assign CALC_SOFTMAX_LOOP_i_mux_rmff = MUX_v_7_2_2(CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_8,
      plm_out_cnsi_wadr_d_reg, or_tmp_337);
  assign CALC_SOFTMAX_LOOP_mux_1_rmff = MUX_v_32_2_2(CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt,
      plm_out_cnsi_d_d_reg, or_tmp_337);
  assign CALC_EXP_LOOP_i_mux_rmff = MUX_v_7_2_2(CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_2,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d_reg,
      or_tmp_339);
  assign ac_math_ac_shift_left_21_1_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_1_rmff
      = MUX_v_67_2_2(operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d_reg,
      or_tmp_339);
  assign or_482_nl = (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1) | exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_4
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0 | (~ COMPUTE_BATCH_LOOP_and_16_tmp)
      | (~ (fsm_output[1]));
  assign CALC_SOFTMAX_LOOP_i_mux_1_rmff = MUX_v_7_2_2(CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_4,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d_reg,
      or_482_nl);
  assign or_483_nl = exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_2 | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1
      | (~ COMPUTE_BATCH_LOOP_and_23_tmp) | (~ (fsm_output[1]));
  assign CALC_EXP_LOOP_i_mux_1_rmff = MUX_v_7_2_2(CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_2_6_0,
      plm_in_cnsi_radr_d_reg, or_483_nl);
  assign softmax_sysc_compute_load_handshake_softmax_sysc_compute_load_handshake_or_rmff
      = (input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_psct & (~(and_dcpl_52
      & (~(CALC_SOFTMAX_LOOP_asn_itm & COMPUTE_BATCH_LOOP_acc_itm_32_1 & COMPUTE_BATCH_LOOP_and_33_tmp))
      & (fsm_output[1])))) | or_tmp_320;
  assign mux_238_nl = MUX_s_1_2_2((~ COMPUTE_BATCH_LOOP_stage_v), nand_tmp_12, COMPUTE_BATCH_LOOP_and_33_tmp);
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_nand_1_cse = ~(mux_238_nl
      & COMPUTE_BATCH_LOOP_stage_0);
  assign CALC_SOFTMAX_LOOP_and_31_cse = compute_wen & (fsm_output[1]);
  assign CALC_SOFTMAX_LOOP_and_72_cse = CALC_SOFTMAX_LOOP_and_31_cse & (~(CALC_SOFTMAX_LOOP_asn_itm
      & (~ COMPUTE_BATCH_LOOP_acc_itm_32_1) & exitL_exit_CALC_SOFTMAX_LOOP_sva))
      & COMPUTE_BATCH_LOOP_and_33_tmp;
  assign and_228_nl = or_107_cse & or_106_cse;
  assign and_227_nl = (plm_out_cns_rls_obj_bawt | (~ CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9)
      | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1) | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0
      | exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9) & or_106_cse;
  assign mux_271_cse = MUX_s_1_2_2(and_228_nl, and_227_nl, plm_out_cnsi_bawt);
  assign nor_95_cse = ~(COMPUTE_BATCH_LOOP_stage_v_8 | (~ mux_tmp_187));
  assign and_232_nl = or_cse & mux_tmp_187;
  assign mux_273_nl = MUX_s_1_2_2(mux_tmp_187, mux_271_cse, reg_COMPUTE_BATCH_LOOP_stage_v_9_cse);
  assign and_231_nl = or_cse & mux_273_nl;
  assign mux_274_nl = MUX_s_1_2_2(and_232_nl, and_231_nl, COMPUTE_BATCH_LOOP_stage_v_7);
  assign mux_275_nl = MUX_s_1_2_2(mux_tmp_187, mux_274_nl, COMPUTE_BATCH_LOOP_stage_v_8);
  assign mux_277_nl = MUX_s_1_2_2(nor_95_cse, mux_275_nl, or_8_cse);
  assign COMPUTE_BATCH_LOOP_and_37_cse = compute_wen & mux_277_nl;
  assign and_826_cse = COMPUTE_BATCH_LOOP_stage_v_7 & COMPUTE_BATCH_LOOP_stage_0_8;
  assign or_8_cse = exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8 | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1)
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0 | CALC_SOFTMAX_LOOP_mul_cmp_bawt;
  assign or_cse = (~ CALC_SOFTMAX_LOOP_asn_itm_8) | exit_COMPUTE_BATCH_LOOP_sva_1_st_8
      | plm_out_cns_req_obj_bawt;
  assign CALC_SOFTMAX_LOOP_and_74_cse = CALC_SOFTMAX_LOOP_and_31_cse & COMPUTE_BATCH_LOOP_and_16_tmp;
  assign CALC_EXP_LOOP_and_5_cse = compute_wen & COMPUTE_BATCH_LOOP_and_19_tmp &
      (fsm_output[1]);
  assign and_837_tmp = ((~ CALC_SOFTMAX_LOOP_asn_1_itm_3) | exit_COMPUTE_BATCH_LOOP_sva_1_3)
      & COMPUTE_BATCH_LOOP_and_19_tmp & (fsm_output[1]);
  assign CALC_EXP_LOOP_i_and_4_cse = COMPUTE_BATCH_LOOP_and_19_tmp & (fsm_output[1]);
  assign COMPUTE_BATCH_LOOP_and_62_cse = CALC_SOFTMAX_LOOP_and_31_cse & COMPUTE_BATCH_LOOP_and_19_tmp;
  assign CALC_SOFTMAX_LOOP_and_75_cse = CALC_SOFTMAX_LOOP_and_31_cse & COMPUTE_BATCH_LOOP_and_23_tmp;
  assign CALC_EXP_LOOP_and_6_cse = CALC_SOFTMAX_LOOP_and_31_cse & COMPUTE_BATCH_LOOP_and_28_tmp;
  assign nor_129_cse = ~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1 | exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_2);
  assign CALC_EXP_LOOP_i_and_3_cse = COMPUTE_BATCH_LOOP_and_28_tmp & (fsm_output[1]);
  assign CALC_SOFTMAX_LOOP_i_and_22_itm = compute_wen & COMPUTE_BATCH_LOOP_and_33_tmp;
  assign and_240_nl = COMPUTE_BATCH_LOOP_stage_0_10 & mux_271_cse;
  assign mux_280_nl = MUX_s_1_2_2(mux_tmp_187, and_240_nl, reg_COMPUTE_BATCH_LOOP_stage_v_9_cse);
  assign and_244_cse = COMPUTE_BATCH_LOOP_stage_0_9 & or_cse & mux_280_nl;
  assign COMPUTE_BATCH_LOOP_and_64_cse = compute_wen & COMPUTE_BATCH_LOOP_and_13_tmp;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_and_cse
      = compute_wen & (~(((~ COMPUTE_BATCH_LOOP_and_16_tmp) & (fsm_output[1])) |
      (fsm_output[0])));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_and_cse = compute_wen
      & COMPUTE_BATCH_LOOP_and_16_tmp & (fsm_output[1]);
  assign COMPUTE_BATCH_LOOP_and_65_cse = compute_wen & COMPUTE_BATCH_LOOP_and_23_tmp
      & (fsm_output[1]);
  assign mux_141_cse = MUX_s_1_2_2((~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1),
      mux_tmp_29, exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign CALC_EXP_LOOP_i_and_2_rgt = and_dcpl_246 & (fsm_output[1]);
  assign nor_127_cse = ~(exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_3 | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1);
  assign CALC_EXP_LOOP_and_7_itm = CALC_SOFTMAX_LOOP_and_31_cse & COMPUTE_BATCH_LOOP_and_33_tmp;
  assign or_106_cse = (~ reg_COMPUTE_BATCH_LOOP_stage_v_10_cse) | output_ready_req_mioi_bawt
      | (~ CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_10) | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_1)
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_0 | exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_10;
  assign or_107_cse = (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1) | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0
      | exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_and_cse = compute_wen
      & (~((~((~ and_dcpl_240) | (~ and_dcpl_220) | (~ and_dcpl_214) | (SUM_EXP_LOOP_acc_1_tmp[73:26]!=48'b000000000000000000000000000000000000000000000000)))
      | or_tmp_20 | (~(CALC_EXP_LOOP_and_svs_st_4 & COMPUTE_BATCH_LOOP_and_16_tmp))
      | (~ (fsm_output[1]))));
  assign CALC_SOFTMAX_LOOP_and_89_cse = CALC_SOFTMAX_LOOP_and_31_cse & (~ exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign COMPUTE_BATCH_LOOP_and_72_cse = compute_wen & COMPUTE_BATCH_LOOP_and_33_tmp
      & (fsm_output[1]);
  assign CALC_SOFTMAX_LOOP_i_and_34_cse = CALC_SOFTMAX_LOOP_and_31_cse & (((~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0)
      & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1 & and_dcpl_246) | and_dcpl_301);
  assign CALC_SOFTMAX_LOOP_i_and_36_cse = CALC_SOFTMAX_LOOP_and_31_cse & (~ or_dcpl_140);
  assign COMPUTE_BATCH_LOOP_stage_0_mx1 = COMPUTE_BATCH_LOOP_stage_0 & (mux_tmp_29
      | (~ exitL_exit_CALC_SOFTMAX_LOOP_sva) | (~ COMPUTE_BATCH_LOOP_and_33_tmp));
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_2_nl = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0
      & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0;
  assign CALC_SOFTMAX_LOOP_mux_24_nl = MUX_s_1_2_2((~ (CALC_SOFTMAX_LOOP_acc_1_tmp[7])),
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1, CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_2_nl);
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1_mx1w0 = (CALC_SOFTMAX_LOOP_mux_24_nl
      & (~ CALC_SOFTMAX_LOOP_and_4_ssc_1)) | CALC_SOFTMAX_LOOP_and_5_ssc_1;
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0_mx1w0 = (lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0
      & (~(CALC_SOFTMAX_LOOP_and_5_ssc_1 | CALC_SOFTMAX_LOOP_equal_tmp_2))) | CALC_SOFTMAX_LOOP_and_4_ssc_1;
  assign exitL_exit_CALC_SOFTMAX_LOOP_sva_mx1w0 = ~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1_mx1w0
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0_mx1w0);
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl
      = MUX_v_10_8_2(10'b1111111101, 10'b1100011001, 10'b1001100100, 10'b0111010000,
      10'b0101010100, 10'b0011101011, 10'b0010010001, 10'b0001000100, operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm[72:70]);
  assign nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm_mx0w1
      = conv_s2u_9_11(ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:10])
      + ({1'b1 , ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl});
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm_mx0w1
      = nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm_mx0w1[10:0];
  assign nl_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm_mx0w1
      = ({1'b1 , (~ libraries_leading_sign_74_0_cfd8a2a1b60025d53198d215150438e7bf24_1)})
      + 8'b00110111;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm_mx0w1
      = nl_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm_mx0w1[7:0];
  assign and_371_nl = and_dcpl_243 & CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_4;
  assign and_372_nl = and_dcpl_243 & (~ CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_4);
  assign or_444_nl = COMPUTE_BATCH_LOOP_asn_2_itm_4 | (~ COMPUTE_BATCH_LOOP_and_16_tmp);
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_mx1
      = MUX1HOT_v_74_3_2(SUM_EXP_LOOP_acc_1_tmp, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_1_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1,
      {and_371_nl , and_372_nl , or_444_nl});
  assign nl_COMPUTE_BATCH_LOOP_acc_nl = ({1'b1 , COMPUTE_BATCH_LOOP_b_sva}) + conv_u2u_32_33(~
      config_batch_sva) + 33'b000000000000000000000000000000001;
  assign COMPUTE_BATCH_LOOP_acc_nl = nl_COMPUTE_BATCH_LOOP_acc_nl[32:0];
  assign COMPUTE_BATCH_LOOP_acc_itm_32_1 = readslicef_33_1_32(COMPUTE_BATCH_LOOP_acc_nl);
  assign nl_SUM_EXP_LOOP_acc_1_tmp = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_1_1
      + conv_u2u_67_74(operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1);
  assign SUM_EXP_LOOP_acc_1_tmp = nl_SUM_EXP_LOOP_acc_1_tmp[73:0];
  assign COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_and_28_nl = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1
      & (~ COMPUTE_BATCH_LOOP_acc_itm_32_1);
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0 = MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1,
      COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_and_28_nl, exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_and_29_nl = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0
      & (~ COMPUTE_BATCH_LOOP_acc_itm_32_1);
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0 = MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0,
      COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_and_29_nl, exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign nl_CALC_SOFTMAX_LOOP_acc_1_tmp = conv_u2u_7_8(CALC_SOFTMAX_LOOP_i_7_0_lpi_1_6_0)
      + 8'b00000001;
  assign CALC_SOFTMAX_LOOP_acc_1_tmp = nl_CALC_SOFTMAX_LOOP_acc_1_tmp[7:0];
  assign COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_11_cse_1 = plm_in_cns_req_obj_bawt
      | (~((~ exit_COMPUTE_BATCH_LOOP_sva_1_st_2) & CALC_SOFTMAX_LOOP_asn_itm_2 &
      COMPUTE_BATCH_LOOP_stage_v_2));
  assign COMPUTE_BATCH_LOOP_or_40_cse_1 = plm_in_cnsi_bawt | (~(nor_127_cse & reg_COMPUTE_BATCH_LOOP_stage_v_3_cse));
  assign COMPUTE_BATCH_LOOP_or_41_cse_1 = plm_in_cns_rls_obj_bawt | (~(CALC_EXP_LOOP_and_svs_st_3
      & CALC_SOFTMAX_LOOP_or_16_cse_1 & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_3)
      & reg_COMPUTE_BATCH_LOOP_stage_v_3_cse));
  assign COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_7_cse_1 = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt
      | (~((~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1 | exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_5))
      & reg_COMPUTE_BATCH_LOOP_stage_v_5_cse));
  assign COMPUTE_BATCH_LOOP_or_4_cse_1 = plm_out_cns_req_obj_bawt | (~((~ exit_COMPUTE_BATCH_LOOP_sva_1_st_8)
      & CALC_SOFTMAX_LOOP_asn_itm_8 & COMPUTE_BATCH_LOOP_stage_v_8));
  assign COMPUTE_BATCH_LOOP_or_10_cse_1 = CALC_SOFTMAX_LOOP_mul_cmp_bawt | (~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0) & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8)
      & COMPUTE_BATCH_LOOP_stage_v_8));
  assign COMPUTE_BATCH_LOOP_or_6_cse_1 = plm_out_cnsi_bawt | (~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0) & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9)
      & reg_COMPUTE_BATCH_LOOP_stage_v_9_cse));
  assign COMPUTE_BATCH_LOOP_or_7_cse_1 = plm_out_cns_rls_obj_bawt | (~(CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9
      & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0)
      & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9) & reg_COMPUTE_BATCH_LOOP_stage_v_9_cse));
  assign COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_1_cse_1 = output_ready_req_mioi_bawt
      | (~(CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_10 & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_1
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_0) & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_10)
      & reg_COMPUTE_BATCH_LOOP_stage_v_10_cse));
  assign CALC_SOFTMAX_LOOP_or_16_cse_1 = (lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1)) | (~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0));
  assign nl_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl
      = $signed((plm_in_cnsi_q_d_mxwt)) * $signed(16'b0101110001010101);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl
      = nl_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl[46:0];
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28
      = readslicef_47_19_28(ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_7_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28[11:10]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_1_nl
      = MUX_v_3_4_2(3'b010, 3'b110, 3'b001, 3'b101, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28[11:10]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = conv_u2u_19_19(({ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_7_nl
      , 1'b0 , ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_1_nl})
      * (ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28[9:0]));
  assign CALC_EXP_LOOP_and_svs_1 = (CALC_EXP_LOOP_acc_1_tmp[7]) & (SUM_EXP_LOOP_acc_2_tmp[7]);
  assign CALC_SOFTMAX_LOOP_or_tmp_1 = (lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0)) | (~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0));
  assign CALC_SOFTMAX_LOOP_equal_tmp_2 = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0);
  assign CALC_SOFTMAX_LOOP_mux_112_nl = MUX_v_7_2_2(CALC_EXP_LOOP_i_7_0_lpi_1_6_0,
      (signext_7_1(~ COMPUTE_BATCH_LOOP_acc_itm_32_1)), exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign nl_CALC_EXP_LOOP_acc_1_tmp = conv_u2u_7_8(CALC_SOFTMAX_LOOP_mux_112_nl)
      + 8'b00000001;
  assign CALC_EXP_LOOP_acc_1_tmp = nl_CALC_EXP_LOOP_acc_1_tmp[7:0];
  assign CALC_SOFTMAX_LOOP_mux_111_nl = MUX_v_7_2_2(SUM_EXP_LOOP_i_7_0_lpi_1_6_0,
      (signext_7_1(~ COMPUTE_BATCH_LOOP_acc_itm_32_1)), exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign nl_SUM_EXP_LOOP_acc_2_tmp = conv_u2u_7_8(CALC_SOFTMAX_LOOP_mux_111_nl) +
      8'b00000001;
  assign SUM_EXP_LOOP_acc_2_tmp = nl_SUM_EXP_LOOP_acc_2_tmp[7:0];
  assign CALC_SOFTMAX_LOOP_and_4_ssc_1 = (~ CALC_EXP_LOOP_and_svs_1) & CALC_SOFTMAX_LOOP_or_tmp_1;
  assign CALC_SOFTMAX_LOOP_and_5_ssc_1 = CALC_EXP_LOOP_and_svs_1 & CALC_SOFTMAX_LOOP_or_tmp_1;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_3_nl
      = MUX_v_8_8_2(8'b00011100, 8'b01001011, 8'b01101100, 8'b10000100, 8'b10010111,
      8'b10100110, 8'b10110011, 8'b10111100, operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm[72:70]);
  assign nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = $signed(({1'b1 , ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_3_nl}))
      * $signed(conv_u2s_10_11(operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm[69:60]));
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:0];
  assign COMPUTE_BATCH_LOOP_and_33_tmp = COMPUTE_BATCH_LOOP_stage_v & (~(COMPUTE_BATCH_LOOP_stage_v_1
      & (~ COMPUTE_BATCH_LOOP_and_28_tmp))) & COMPUTE_BATCH_LOOP_stage_0_1 & COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_11_cse_1
      & COMPUTE_BATCH_LOOP_or_40_cse_1 & COMPUTE_BATCH_LOOP_or_41_cse_1 & COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_7_cse_1
      & COMPUTE_BATCH_LOOP_or_4_cse_1 & COMPUTE_BATCH_LOOP_or_10_cse_1 & COMPUTE_BATCH_LOOP_or_6_cse_1
      & COMPUTE_BATCH_LOOP_or_7_cse_1 & COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_1_cse_1;
  assign COMPUTE_BATCH_LOOP_and_28_tmp = COMPUTE_BATCH_LOOP_stage_v_1 & (~(COMPUTE_BATCH_LOOP_stage_v_2
      & (~ COMPUTE_BATCH_LOOP_and_23_tmp))) & COMPUTE_BATCH_LOOP_stage_0_2 & (input_ready_ack_mioi_bawt
      | (~((~ exit_COMPUTE_BATCH_LOOP_sva_1_st_1) & CALC_SOFTMAX_LOOP_asn_itm_1)))
      & COMPUTE_BATCH_LOOP_or_40_cse_1 & COMPUTE_BATCH_LOOP_or_41_cse_1 & COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_7_cse_1
      & COMPUTE_BATCH_LOOP_or_4_cse_1 & COMPUTE_BATCH_LOOP_or_10_cse_1 & COMPUTE_BATCH_LOOP_or_6_cse_1
      & COMPUTE_BATCH_LOOP_or_7_cse_1 & COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_1_cse_1;
  assign COMPUTE_BATCH_LOOP_and_23_tmp = COMPUTE_BATCH_LOOP_stage_v_2 & (~(reg_COMPUTE_BATCH_LOOP_stage_v_3_cse
      & (~ COMPUTE_BATCH_LOOP_and_19_tmp))) & COMPUTE_BATCH_LOOP_stage_0_3 & COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_11_cse_1
      & COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_7_cse_1 & COMPUTE_BATCH_LOOP_or_4_cse_1
      & COMPUTE_BATCH_LOOP_or_10_cse_1 & COMPUTE_BATCH_LOOP_or_6_cse_1 & COMPUTE_BATCH_LOOP_or_7_cse_1
      & COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_1_cse_1;
  assign COMPUTE_BATCH_LOOP_and_19_tmp = reg_COMPUTE_BATCH_LOOP_stage_v_3_cse & (~(COMPUTE_BATCH_LOOP_stage_v_4
      & (~ COMPUTE_BATCH_LOOP_and_16_tmp))) & COMPUTE_BATCH_LOOP_stage_0_4 & (plm_in_cnsi_bawt
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1 | exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_3)
      & (plm_in_cns_rls_obj_bawt | (~(CALC_EXP_LOOP_and_svs_st_3 & CALC_SOFTMAX_LOOP_or_16_cse_1
      & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_3)))) & COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_7_cse_1
      & COMPUTE_BATCH_LOOP_or_4_cse_1 & COMPUTE_BATCH_LOOP_or_10_cse_1 & COMPUTE_BATCH_LOOP_or_6_cse_1
      & COMPUTE_BATCH_LOOP_or_7_cse_1 & COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_1_cse_1;
  assign COMPUTE_BATCH_LOOP_and_16_tmp = COMPUTE_BATCH_LOOP_stage_v_4 & (~(reg_COMPUTE_BATCH_LOOP_stage_v_5_cse
      & (~ COMPUTE_BATCH_LOOP_and_13_tmp))) & COMPUTE_BATCH_LOOP_stage_0_5 & COMPUTE_BATCH_LOOP_or_4_cse_1
      & COMPUTE_BATCH_LOOP_or_10_cse_1 & COMPUTE_BATCH_LOOP_or_6_cse_1 & COMPUTE_BATCH_LOOP_or_7_cse_1
      & COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_1_cse_1;
  assign or_634_nl = COMPUTE_BATCH_LOOP_stage_v_8 | mux_248_cse;
  assign nand_23_nl = ~(COMPUTE_BATCH_LOOP_stage_0_8 & mux_244_cse);
  assign mux_256_nl = MUX_s_1_2_2(or_tmp_202, nand_23_nl, or_cse);
  assign mux_258_nl = MUX_s_1_2_2((~ mux_tmp_229), mux_256_nl, COMPUTE_BATCH_LOOP_stage_v_7);
  assign mux_260_nl = MUX_s_1_2_2(or_634_nl, mux_258_nl, or_8_cse);
  assign COMPUTE_BATCH_LOOP_and_13_tmp = reg_COMPUTE_BATCH_LOOP_stage_v_5_cse & (~(COMPUTE_BATCH_LOOP_stage_v_6
      & (mux_260_nl | or_dcpl_50))) & COMPUTE_BATCH_LOOP_stage_0_6 & (ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1 | exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_5)
      & COMPUTE_BATCH_LOOP_or_4_cse_1 & COMPUTE_BATCH_LOOP_or_10_cse_1 & COMPUTE_BATCH_LOOP_or_6_cse_1
      & COMPUTE_BATCH_LOOP_or_7_cse_1 & COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_or_1_cse_1;
  assign and_23_cse = or_181_cse & plm_out_cnsi_bawt & or_106_cse;
  assign nor_1_nl = ~((~ reg_COMPUTE_BATCH_LOOP_stage_v_9_cse) | exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0 | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1));
  assign mux_tmp_1 = MUX_s_1_2_2(or_106_cse, and_23_cse, nor_1_nl);
  assign nor_3_cse = ~(exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9 | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0
      | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1));
  assign mux_21_cse = MUX_s_1_2_2(or_106_cse, and_23_cse, nor_3_cse);
  assign or_tmp_20 = exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_4 | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1;
  assign mux_tmp_29 = MUX_s_1_2_2((~ CALC_SOFTMAX_LOOP_asn_itm), CALC_SOFTMAX_LOOP_asn_itm,
      COMPUTE_BATCH_LOOP_acc_itm_32_1);
  assign nor_tmp_12 = COMPUTE_BATCH_LOOP_stage_v_6 & COMPUTE_BATCH_LOOP_stage_0_7;
  assign or_48_cse = (~ reg_COMPUTE_BATCH_LOOP_stage_v_9_cse) | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1)
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0 | exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9;
  assign or_46_cse = plm_out_cns_rls_obj_bawt | (~ CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9)
      | (~ reg_COMPUTE_BATCH_LOOP_stage_v_9_cse) | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1)
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0 | exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9;
  assign or_120_cse = output_ready_req_mioi_bawt | (~ CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_10)
      | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_1) | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_0
      | exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_10;
  assign and_dcpl_52 = CALC_SOFTMAX_LOOP_asn_itm_1 & COMPUTE_BATCH_LOOP_and_28_tmp
      & (~ exit_COMPUTE_BATCH_LOOP_sva_1_st_1);
  assign and_dcpl_54 = CALC_SOFTMAX_LOOP_asn_itm_2 & COMPUTE_BATCH_LOOP_and_23_tmp
      & (~ exit_COMPUTE_BATCH_LOOP_sva_1_st_2);
  assign and_111_nl = or_48_cse & or_106_cse;
  assign and_110_nl = or_46_cse & or_106_cse;
  assign mux_tmp_187 = MUX_s_1_2_2(and_111_nl, and_110_nl, plm_out_cnsi_bawt);
  assign mux_206_nl = MUX_s_1_2_2(mux_tmp_187, and_244_cse, COMPUTE_BATCH_LOOP_stage_v_8);
  assign mux_tmp_190 = MUX_s_1_2_2(nor_95_cse, mux_206_nl, or_8_cse);
  assign and_dcpl_64 = COMPUTE_BATCH_LOOP_stage_0_9 & plm_out_cns_req_obj_bawt &
      (~ exit_COMPUTE_BATCH_LOOP_sva_1_st_8) & CALC_SOFTMAX_LOOP_asn_itm_8 & COMPUTE_BATCH_LOOP_stage_v_8;
  assign and_119_nl = COMPUTE_BATCH_LOOP_stage_0_10 & or_106_cse;
  assign mux_tmp_191 = MUX_s_1_2_2(or_106_cse, and_119_nl, reg_COMPUTE_BATCH_LOOP_stage_v_9_cse);
  assign or_tmp_152 = reg_COMPUTE_BATCH_LOOP_stage_v_9_cse | (~ or_106_cse);
  assign mux_209_nl = MUX_s_1_2_2(mux_tmp_191, (~ or_tmp_152), CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9);
  assign mux_210_nl = MUX_s_1_2_2(mux_209_nl, mux_tmp_191, plm_out_cns_rls_obj_bawt);
  assign mux_211_nl = MUX_s_1_2_2((~ or_tmp_152), mux_210_nl, plm_out_cnsi_bawt);
  assign mux_212_cse = MUX_s_1_2_2(mux_211_nl, mux_tmp_191, or_107_cse);
  assign and_dcpl_82 = (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_0) & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_1
      & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_10) & CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_10
      & output_ready_req_mioi_bawt & reg_COMPUTE_BATCH_LOOP_stage_v_10_cse;
  assign and_dcpl_84 = (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9) & reg_COMPUTE_BATCH_LOOP_stage_v_9_cse
      & COMPUTE_BATCH_LOOP_stage_0_10;
  assign and_dcpl_103 = COMPUTE_BATCH_LOOP_stage_0_9 & CALC_SOFTMAX_LOOP_mul_cmp_bawt;
  assign and_dcpl_106 = mux_212_cse & or_cse;
  assign and_tmp_54 = or_8_cse & mux_212_cse;
  assign or_dcpl_16 = ~(reg_COMPUTE_BATCH_LOOP_stage_v_9_cse & COMPUTE_BATCH_LOOP_stage_0_10);
  assign and_dcpl_121 = (~(plm_out_cns_req_obj_bawt | exit_COMPUTE_BATCH_LOOP_sva_1_st_8))
      & CALC_SOFTMAX_LOOP_asn_itm_8;
  assign nand_tmp_12 = ~(exitL_exit_CALC_SOFTMAX_LOOP_sva & (~ mux_tmp_29));
  assign and_dcpl_125 = (~ mux_tmp_29) & exitL_exit_CALC_SOFTMAX_LOOP_sva;
  assign or_dcpl_45 = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0 | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1);
  assign or_tmp_202 = (~ COMPUTE_BATCH_LOOP_stage_0_8) | COMPUTE_BATCH_LOOP_stage_v_8
      | (~ mux_tmp_187);
  assign mux_tmp_229 = MUX_s_1_2_2(nor_95_cse, mux_tmp_187, or_cse);
  assign mux_241_nl = MUX_s_1_2_2(mux_tmp_187, mux_271_cse, COMPUTE_BATCH_LOOP_stage_v_8);
  assign mux_242_nl = MUX_s_1_2_2(nor_95_cse, mux_241_nl, COMPUTE_BATCH_LOOP_stage_0_10);
  assign mux_243_cse = MUX_s_1_2_2(mux_tmp_187, mux_242_nl, reg_COMPUTE_BATCH_LOOP_stage_v_9_cse);
  assign mux_244_cse = MUX_s_1_2_2(nor_95_cse, mux_243_cse, COMPUTE_BATCH_LOOP_stage_0_9);
  assign mux_248_cse = MUX_s_1_2_2((~ mux_tmp_229), or_tmp_202, COMPUTE_BATCH_LOOP_stage_v_7);
  assign nor_98_nl = ~(COMPUTE_BATCH_LOOP_stage_v_8 | mux_248_cse);
  assign and_210_nl = COMPUTE_BATCH_LOOP_stage_0_8 & mux_244_cse;
  assign mux_245_nl = MUX_s_1_2_2((~ or_tmp_202), and_210_nl, or_cse);
  assign mux_247_nl = MUX_s_1_2_2(mux_tmp_229, mux_245_nl, COMPUTE_BATCH_LOOP_stage_v_7);
  assign mux_tmp_232 = MUX_s_1_2_2(nor_98_nl, mux_247_nl, or_8_cse);
  assign or_dcpl_50 = ~(COMPUTE_BATCH_LOOP_stage_v_6 & COMPUTE_BATCH_LOOP_stage_0_7);
  assign and_dcpl_140 = mux_tmp_232 & nor_tmp_12;
  assign and_226_cse = nor_tmp_12 & mux_tmp_229;
  assign or_dcpl_52 = ~(COMPUTE_BATCH_LOOP_stage_0_8 & COMPUTE_BATCH_LOOP_stage_v_7);
  assign and_dcpl_142 = COMPUTE_BATCH_LOOP_stage_0_9 & COMPUTE_BATCH_LOOP_stage_v_8;
  assign and_dcpl_144 = and_tmp_54 & or_cse;
  assign and_tmp_85 = COMPUTE_BATCH_LOOP_stage_v_7 & COMPUTE_BATCH_LOOP_stage_0_8
      & mux_tmp_187;
  assign or_dcpl_53 = (~ mux_tmp_190) | or_dcpl_52;
  assign mux_22_nl = MUX_s_1_2_2(mux_tmp_1, mux_21_cse, reg_COMPUTE_BATCH_LOOP_stage_v_9_cse);
  assign and_256_nl = or_8_cse & or_cse & mux_22_nl;
  assign mux_291_itm = MUX_s_1_2_2(mux_tmp_1, and_256_nl, COMPUTE_BATCH_LOOP_stage_v_8);
  assign and_dcpl_147 = reg_COMPUTE_BATCH_LOOP_stage_v_9_cse & COMPUTE_BATCH_LOOP_stage_0_10;
  assign or_dcpl_56 = (~(or_8_cse & mux_212_cse)) | and_dcpl_121 | (~ COMPUTE_BATCH_LOOP_stage_0_9)
      | (~ COMPUTE_BATCH_LOOP_stage_v_8);
  assign or_dcpl_57 = (~ mux_21_cse) | or_dcpl_16;
  assign and_dcpl_165 = exitL_exit_CALC_SOFTMAX_LOOP_sva & COMPUTE_BATCH_LOOP_and_33_tmp;
  assign and_dcpl_166 = (~ mux_tmp_29) & and_dcpl_165;
  assign and_dcpl_214 = ~((SUM_EXP_LOOP_acc_1_tmp[25:24]!=2'b00));
  assign and_dcpl_220 = (SUM_EXP_LOOP_acc_1_tmp[23:19]==5'b00000);
  assign and_dcpl_240 = (SUM_EXP_LOOP_acc_1_tmp[18:0]==19'b0000000000000000000);
  assign and_dcpl_243 = (~ COMPUTE_BATCH_LOOP_asn_2_itm_4) & COMPUTE_BATCH_LOOP_and_16_tmp;
  assign and_dcpl_246 = (~ exitL_exit_CALC_SOFTMAX_LOOP_sva) & COMPUTE_BATCH_LOOP_and_33_tmp;
  assign or_dcpl_140 = or_dcpl_45 | exitL_exit_CALC_SOFTMAX_LOOP_sva;
  assign and_dcpl_301 = or_dcpl_140 & COMPUTE_BATCH_LOOP_and_33_tmp;
  assign or_tmp_309 = and_dcpl_52 & (fsm_output[1]);
  assign or_tmp_320 = CALC_SOFTMAX_LOOP_asn_itm & COMPUTE_BATCH_LOOP_acc_itm_32_1
      & COMPUTE_BATCH_LOOP_and_33_tmp & (fsm_output[1]);
  assign or_tmp_322 = or_106_cse & plm_out_cnsi_bawt & plm_out_cns_rls_obj_bawt &
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9 & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0) & and_dcpl_84 & (fsm_output[1]);
  assign or_tmp_337 = (~ mux_212_cse) | and_dcpl_121 | (~ COMPUTE_BATCH_LOOP_stage_0_9)
      | (~ CALC_SOFTMAX_LOOP_mul_cmp_bawt) | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0
      | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1) | exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8
      | (~ COMPUTE_BATCH_LOOP_stage_v_8) | (~ (fsm_output[1]));
  assign or_tmp_339 = or_tmp_20 | (~ COMPUTE_BATCH_LOOP_and_16_tmp) | (~ (fsm_output[1]));
  assign or_tmp_431 = ~((~ and_dcpl_240) | (~ and_dcpl_220) | (~ and_dcpl_214) |
      (SUM_EXP_LOOP_acc_1_tmp[73:26]!=48'b000000000000000000000000000000000000000000000000)
      | (~ COMPUTE_BATCH_LOOP_and_16_tmp) | (~ (fsm_output[1])));
  assign plm_in_cns_req_obj_iswt0_mx0c1 = and_dcpl_54 & ((~(CALC_SOFTMAX_LOOP_asn_itm_1
      & COMPUTE_BATCH_LOOP_and_28_tmp)) | exit_COMPUTE_BATCH_LOOP_sva_1_st_1) & (fsm_output[1]);
  assign nor_78_nl = ~(COMPUTE_BATCH_LOOP_stage_0_8 | (~ mux_212_cse));
  assign or_154_nl = (~ COMPUTE_BATCH_LOOP_stage_v_7) | (~ CALC_SOFTMAX_LOOP_asn_itm_7)
      | exit_COMPUTE_BATCH_LOOP_sva_1_st_7;
  assign mux_213_nl = MUX_s_1_2_2(nor_78_nl, mux_212_cse, or_154_nl);
  assign plm_out_cns_req_obj_iswt0_mx0c1 = or_8_cse & mux_213_nl & and_dcpl_64 &
      (fsm_output[1]);
  assign COMPUTE_BATCH_LOOP_stage_v_6_mx0c1 = COMPUTE_BATCH_LOOP_and_13_tmp & (fsm_output[1]);
  assign COMPUTE_BATCH_LOOP_stage_v_7_mx0c1 = and_dcpl_140 & (fsm_output[1]);
  assign COMPUTE_BATCH_LOOP_stage_0_7_mx0c1 = (and_dcpl_140 | COMPUTE_BATCH_LOOP_and_13_tmp)
      & (fsm_output[1]);
  assign mux_269_nl = MUX_s_1_2_2((~ and_226_cse), or_tmp_202, COMPUTE_BATCH_LOOP_stage_v_7);
  assign nor_106_nl = ~(COMPUTE_BATCH_LOOP_stage_v_8 | mux_269_nl);
  assign and_813_nl = or_cse & COMPUTE_BATCH_LOOP_stage_0_9;
  assign mux_266_nl = MUX_s_1_2_2(nor_95_cse, mux_243_cse, and_813_nl);
  assign and_225_nl = COMPUTE_BATCH_LOOP_stage_0_8 & mux_266_nl;
  assign mux_268_nl = MUX_s_1_2_2(and_226_cse, and_225_nl, COMPUTE_BATCH_LOOP_stage_v_7);
  assign mux_270_nl = MUX_s_1_2_2(nor_106_nl, mux_268_nl, or_8_cse);
  assign COMPUTE_BATCH_LOOP_stage_0_8_mx0c1 = mux_270_nl & (fsm_output[1]);
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d
      = ac_math_ac_shift_left_21_1_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_1_rmff;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d
      = CALC_SOFTMAX_LOOP_i_mux_1_rmff;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d
      = CALC_EXP_LOOP_i_mux_rmff;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  assign plm_in_cnsi_radr_d = CALC_EXP_LOOP_i_mux_1_rmff;
  assign plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d = plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_reg;
  assign plm_out_cnsi_d_d = CALC_SOFTMAX_LOOP_mux_1_rmff;
  assign plm_out_cnsi_wadr_d = CALC_SOFTMAX_LOOP_i_mux_rmff;
  assign plm_out_cnsi_we_d_pff = plm_out_cnsi_we_d_iff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cns_req_obj_iswt0 <= 1'b0;
    end
    else if ( compute_wen & (or_tmp_309 | plm_in_cns_req_obj_iswt0_mx0c1) ) begin
      plm_in_cns_req_obj_iswt0 <= ~ plm_in_cns_req_obj_iswt0_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cns_req_obj_iswt0 <= 1'b0;
    end
    else if ( compute_wen & ((mux_tmp_190 & and_826_cse & CALC_SOFTMAX_LOOP_asn_itm_7
        & (~ exit_COMPUTE_BATCH_LOOP_sva_1_st_7) & (fsm_output[1])) | plm_out_cns_req_obj_iswt0_mx0c1)
        ) begin
      plm_out_cns_req_obj_iswt0 <= ~ plm_out_cns_req_obj_iswt0_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( compute_wen ) begin
      output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_psct <= softmax_sysc_compute_store_handshake_softmax_sysc_compute_store_handshake_or_rmff;
      plm_out_cnsi_wadr_d_reg <= CALC_SOFTMAX_LOOP_i_mux_rmff;
      plm_out_cnsi_d_d_reg <= CALC_SOFTMAX_LOOP_mux_1_rmff;
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d_reg
          <= CALC_EXP_LOOP_i_mux_rmff;
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d_reg
          <= ac_math_ac_shift_left_21_1_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_1_rmff;
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d_reg
          <= CALC_SOFTMAX_LOOP_i_mux_1_rmff;
      plm_in_cnsi_radr_d_reg <= CALC_EXP_LOOP_i_mux_1_rmff;
      input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_psct <= softmax_sysc_compute_load_handshake_softmax_sysc_compute_load_handshake_or_rmff;
      COMPUTE_BATCH_LOOP_b_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          COMPUTE_BATCH_LOOP_b_mux_nl, (fsm_output[1]));
      config_batch_sva <= MUX_v_32_2_2(conf_info, config_batch_sva, fsm_output[1]);
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_8 <= MUX_v_7_2_2(CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_8,
          CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_7, mux_291_itm);
      reg_COMPUTE_BATCH_LOOP_stage_v_5_cse <= ((reg_COMPUTE_BATCH_LOOP_stage_v_5_cse
          & (~ COMPUTE_BATCH_LOOP_and_13_tmp)) | COMPUTE_BATCH_LOOP_and_16_tmp) &
          (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_v_4 <= ((COMPUTE_BATCH_LOOP_stage_v_4 & (~ COMPUTE_BATCH_LOOP_and_16_tmp))
          | COMPUTE_BATCH_LOOP_and_19_tmp) & (fsm_output[1]);
      CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_2 <= MUX_v_7_2_2(CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_2,
          CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_1, CALC_EXP_LOOP_i_and_4_cse);
      ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_itm_1
          <= MUX_v_11_2_2(ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_itm_1,
          ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl,
          CALC_EXP_LOOP_i_and_4_cse);
      ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18_0_1_itm_1
          <= MUX_v_10_2_2(ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_sdt_18_0_1_itm_1,
          (ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[9:0]),
          CALC_EXP_LOOP_i_and_4_cse);
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_32_14_18_12_itm_1
          <= MUX_v_7_2_2(ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_32_14_18_12_itm_1,
          (ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28[18:12]),
          CALC_EXP_LOOP_i_and_4_cse);
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_4 <= MUX_v_7_2_2(CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_4,
          CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_3, CALC_EXP_LOOP_i_and_4_cse);
      reg_COMPUTE_BATCH_LOOP_stage_v_3_cse <= ((reg_COMPUTE_BATCH_LOOP_stage_v_3_cse
          & (~ COMPUTE_BATCH_LOOP_and_19_tmp)) | COMPUTE_BATCH_LOOP_and_23_tmp) &
          (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_v_2 <= ((COMPUTE_BATCH_LOOP_stage_v_2 & (~ COMPUTE_BATCH_LOOP_and_23_tmp))
          | COMPUTE_BATCH_LOOP_and_28_tmp) & (fsm_output[1]);
      CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_2_6_0 <= MUX_v_7_2_2(CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_2_6_0,
          CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_1_6_0, CALC_EXP_LOOP_i_and_3_cse);
      COMPUTE_BATCH_LOOP_stage_v_1 <= ((COMPUTE_BATCH_LOOP_stage_v_1 & (~ COMPUTE_BATCH_LOOP_and_28_tmp))
          | COMPUTE_BATCH_LOOP_and_33_tmp) & (fsm_output[1]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_cse
          <= 1'b0;
      reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_1_cse
          <= 1'b0;
      reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_cse
          <= 1'b0;
      input_ready_ack_mioi_iswt0 <= 1'b0;
      reg_output_ready_req_mioi_iswt0_cse <= 1'b0;
      reg_plm_in_cnsi_iswt0_cse <= 1'b0;
      reg_plm_out_cnsi_iswt0_cse <= 1'b0;
      reg_plm_out_cns_rls_obj_iswt0_cse <= 1'b0;
      reg_plm_in_cns_rls_obj_iswt0_cse <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_v <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm <= 1'b0;
      exitL_exit_CALC_SOFTMAX_LOOP_sva <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_v_8 <= 1'b0;
      reg_COMPUTE_BATCH_LOOP_stage_v_9_cse <= 1'b0;
      reg_COMPUTE_BATCH_LOOP_stage_v_10_cse <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_1 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_2 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_3 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_4 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_5 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_6 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_9 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_10 <= 1'b0;
    end
    else if ( compute_wen ) begin
      reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_cse
          <= and_443_rmff;
      reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_1_cse
          <= and_445_rmff;
      reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_cse
          <= and_447_rmff;
      input_ready_ack_mioi_iswt0 <= or_tmp_320;
      reg_output_ready_req_mioi_iswt0_cse <= or_tmp_322;
      reg_plm_in_cnsi_iswt0_cse <= and_459_rmff;
      reg_plm_out_cnsi_iswt0_cse <= and_463_rmff;
      reg_plm_out_cns_rls_obj_iswt0_cse <= and_dcpl_106 & and_dcpl_103 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0)
          & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1 & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8)
          & COMPUTE_BATCH_LOOP_stage_v_8 & CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_8
          & (fsm_output[1]);
      reg_plm_in_cns_rls_obj_iswt0_cse <= nor_129_cse & COMPUTE_BATCH_LOOP_and_23_tmp
          & CALC_EXP_LOOP_and_svs_st_2 & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_v <= ~((~(COMPUTE_BATCH_LOOP_stage_v & (~((and_dcpl_125
          | (~ COMPUTE_BATCH_LOOP_stage_0)) & COMPUTE_BATCH_LOOP_and_33_tmp)))) &
          ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_nand_1_cse &
          (fsm_output[1]));
      COMPUTE_BATCH_LOOP_stage_0 <= COMPUTE_BATCH_LOOP_stage_0_mx1 | (~ (fsm_output[1]));
      CALC_SOFTMAX_LOOP_asn_itm <= COMPUTE_BATCH_LOOP_mux1h_nl | (~ (fsm_output[1]));
      exitL_exit_CALC_SOFTMAX_LOOP_sva <= COMPUTE_BATCH_LOOP_mux_86_nl | (~ (fsm_output[1]));
      COMPUTE_BATCH_LOOP_stage_v_8 <= ((COMPUTE_BATCH_LOOP_stage_v_8 & (~(and_dcpl_144
          & and_dcpl_142 & or_dcpl_52))) | (mux_tmp_190 & and_826_cse)) & (fsm_output[1]);
      reg_COMPUTE_BATCH_LOOP_stage_v_9_cse <= ((reg_COMPUTE_BATCH_LOOP_stage_v_9_cse
          & (~(mux_293_nl & and_dcpl_147))) | (and_dcpl_144 & and_dcpl_142)) & (fsm_output[1]);
      reg_COMPUTE_BATCH_LOOP_stage_v_10_cse <= ((reg_COMPUTE_BATCH_LOOP_stage_v_10_cse
          & (~ mux_302_nl)) | (mux_21_cse & and_dcpl_147)) & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_1 <= ~((~(operator_74_54_false_AC_TRN_AC_WRAP_1_mux_nl
          & (~ and_dcpl_166))) & (fsm_output[1]));
      COMPUTE_BATCH_LOOP_stage_0_2 <= COMPUTE_BATCH_LOOP_mux_85_nl & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_3 <= COMPUTE_BATCH_LOOP_mux_84_nl & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_4 <= COMPUTE_BATCH_LOOP_mux_83_nl & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_5 <= COMPUTE_BATCH_LOOP_mux_82_nl & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_6 <= COMPUTE_BATCH_LOOP_mux_81_nl & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_9 <= COMPUTE_BATCH_LOOP_mux_80_nl & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_10 <= COMPUTE_BATCH_LOOP_mux_79_nl & (fsm_output[1]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0 <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_72_cse ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1_mx1w0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0_mx1w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      COMPUTE_BATCH_LOOP_stage_v_6 <= 1'b0;
    end
    else if ( compute_wen & ((mux_tmp_232 & nor_tmp_12 & (~ COMPUTE_BATCH_LOOP_and_13_tmp)
        & (fsm_output[1])) | (fsm_output[0]) | COMPUTE_BATCH_LOOP_stage_v_6_mx0c1)
        ) begin
      COMPUTE_BATCH_LOOP_stage_v_6 <= COMPUTE_BATCH_LOOP_stage_v_6_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      COMPUTE_BATCH_LOOP_stage_v_7 <= 1'b0;
    end
    else if ( compute_wen & ((mux_tmp_190 & and_826_cse & or_dcpl_50 & (fsm_output[1]))
        | (fsm_output[0]) | COMPUTE_BATCH_LOOP_stage_v_7_mx0c1) ) begin
      COMPUTE_BATCH_LOOP_stage_v_7 <= COMPUTE_BATCH_LOOP_stage_v_7_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( COMPUTE_BATCH_LOOP_and_37_cse ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_7 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_COMPUTE_BATCH_LOOP_sva_1_st_7 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_7 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_7 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_7 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0 <= 1'b0;
    end
    else if ( COMPUTE_BATCH_LOOP_and_37_cse ) begin
      exit_COMPUTE_BATCH_LOOP_sva_1_st_7 <= exit_COMPUTE_BATCH_LOOP_sva_1_st_6;
      CALC_SOFTMAX_LOOP_asn_itm_7 <= CALC_SOFTMAX_LOOP_asn_itm_6;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_7 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_6;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_7 <= exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_6;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0;
    end
  end
  always @(posedge clk) begin
    if ( CALC_SOFTMAX_LOOP_and_31_cse ) begin
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1
          <= ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_mx1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_COMPUTE_BATCH_LOOP_sva_1_st_8 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_8 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_10 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_0 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_10 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_5 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_4 <= 1'b0;
      CALC_EXP_LOOP_and_svs_st_3 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_3 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_2 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_2 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_1 <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_31_cse ) begin
      exit_COMPUTE_BATCH_LOOP_sva_1_st_8 <= MUX_s_1_2_2(exit_COMPUTE_BATCH_LOOP_sva_1_st_7,
          exit_COMPUTE_BATCH_LOOP_sva_1_st_8, or_dcpl_53);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1, or_dcpl_53);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0, or_dcpl_53);
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8 <= MUX_s_1_2_2(exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_7,
          exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8, or_dcpl_53);
      CALC_SOFTMAX_LOOP_asn_itm_8 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_asn_itm_7, CALC_SOFTMAX_LOOP_asn_itm_8,
          or_dcpl_53);
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_8,
          CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9, or_dcpl_56);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1, or_dcpl_56);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0, or_dcpl_56);
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9 <= MUX_s_1_2_2(exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8,
          exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9, or_dcpl_56);
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_10 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9,
          CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_10, or_dcpl_57);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_1, or_dcpl_57);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_0 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_10_0, or_dcpl_57);
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_10 <= MUX_s_1_2_2(exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9,
          exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_10, or_dcpl_57);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1, COMPUTE_BATCH_LOOP_and_16_tmp);
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_5 <= MUX_s_1_2_2(exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_5,
          exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_4, COMPUTE_BATCH_LOOP_and_16_tmp);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1, COMPUTE_BATCH_LOOP_and_19_tmp);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0, COMPUTE_BATCH_LOOP_and_19_tmp);
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_4 <= MUX_s_1_2_2(exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_4,
          exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_3, COMPUTE_BATCH_LOOP_and_19_tmp);
      CALC_EXP_LOOP_and_svs_st_3 <= MUX_s_1_2_2(CALC_EXP_LOOP_and_svs_st_3, CALC_EXP_LOOP_and_svs_st_2,
          COMPUTE_BATCH_LOOP_and_23_tmp);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1, COMPUTE_BATCH_LOOP_and_23_tmp);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0, COMPUTE_BATCH_LOOP_and_23_tmp);
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_3 <= MUX_s_1_2_2(exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_3,
          exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_2, COMPUTE_BATCH_LOOP_and_23_tmp);
      exit_COMPUTE_BATCH_LOOP_sva_1_st_2 <= MUX_s_1_2_2(exit_COMPUTE_BATCH_LOOP_sva_1_st_2,
          exit_COMPUTE_BATCH_LOOP_sva_1_st_1, COMPUTE_BATCH_LOOP_and_28_tmp);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1, COMPUTE_BATCH_LOOP_and_28_tmp);
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_2 <= MUX_s_1_2_2(exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_2,
          exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_1, COMPUTE_BATCH_LOOP_and_28_tmp);
      CALC_SOFTMAX_LOOP_asn_itm_2 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_asn_itm_2, CALC_SOFTMAX_LOOP_asn_itm_1,
          COMPUTE_BATCH_LOOP_and_28_tmp);
      exit_COMPUTE_BATCH_LOOP_sva_1_st_1 <= MUX1HOT_s_1_3_2((~ COMPUTE_BATCH_LOOP_acc_itm_32_1),
          exit_COMPUTE_BATCH_LOOP_sva_1_st, exit_COMPUTE_BATCH_LOOP_sva_1_st_1, {and_284_nl
          , and_285_nl , (~ COMPUTE_BATCH_LOOP_and_33_tmp)});
      CALC_SOFTMAX_LOOP_asn_itm_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_asn_itm_1, CALC_SOFTMAX_LOOP_asn_itm,
          COMPUTE_BATCH_LOOP_and_33_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_8 <= 1'b0;
    end
    else if ( compute_wen & mux_291_itm ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_8 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( compute_wen & (~ COMPUTE_BATCH_LOOP_asn_2_itm_5) & CALC_SOFTMAX_LOOP_and_10_itm_5
        & COMPUTE_BATCH_LOOP_and_13_tmp & (fsm_output[1]) ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1
          <= MUX_v_94_2_2(operator_94_21_false_AC_TRN_AC_WRAP_rshift_itm, 94'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
          ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_itm_1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_0 <= 1'b0;
      COMPUTE_BATCH_LOOP_asn_2_itm_5 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_5 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_5 <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_74_cse ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0;
      COMPUTE_BATCH_LOOP_asn_2_itm_5 <= COMPUTE_BATCH_LOOP_asn_2_itm_4;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_5 <= exit_COMPUTE_BATCH_LOOP_sva_1_st_4;
      CALC_SOFTMAX_LOOP_asn_itm_5 <= CALC_SOFTMAX_LOOP_asn_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_EXP_LOOP_and_svs_st_4 <= 1'b0;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_4 <= 1'b0;
    end
    else if ( CALC_EXP_LOOP_and_5_cse ) begin
      CALC_EXP_LOOP_and_svs_st_4 <= CALC_EXP_LOOP_and_svs_st_3;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_4 <= CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( compute_wen & ((CALC_SOFTMAX_LOOP_asn_1_itm_3 & COMPUTE_BATCH_LOOP_and_19_tmp
        & (fsm_output[1])) | and_837_tmp) ) begin
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_1_1
          <= MUX_v_74_2_2(({{73{exit_COMPUTE_BATCH_LOOP_sva_1_3}}, exit_COMPUTE_BATCH_LOOP_sva_1_3}),
          ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_mx1,
          and_837_tmp);
    end
  end
  always @(posedge clk) begin
    if ( COMPUTE_BATCH_LOOP_and_62_cse ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_4 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      COMPUTE_BATCH_LOOP_asn_2_itm_4 <= 1'b0;
      CALC_SOFTMAX_LOOP_and_10_itm_4 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_4 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_4 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_4 <= 1'b0;
    end
    else if ( COMPUTE_BATCH_LOOP_and_62_cse ) begin
      COMPUTE_BATCH_LOOP_asn_2_itm_4 <= COMPUTE_BATCH_LOOP_asn_2_itm_3;
      CALC_SOFTMAX_LOOP_and_10_itm_4 <= CALC_SOFTMAX_LOOP_and_10_itm_3;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_4 <= exit_COMPUTE_BATCH_LOOP_sva_1_st_3;
      CALC_SOFTMAX_LOOP_asn_itm_4 <= CALC_SOFTMAX_LOOP_asn_itm_3;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_4 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( CALC_SOFTMAX_LOOP_and_75_cse ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_3 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_asn_itm_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_1_itm_3 <= 1'b0;
      COMPUTE_BATCH_LOOP_asn_2_itm_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_and_10_itm_3 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_3 <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_75_cse ) begin
      CALC_SOFTMAX_LOOP_asn_itm_3 <= CALC_SOFTMAX_LOOP_asn_itm_2;
      CALC_SOFTMAX_LOOP_asn_1_itm_3 <= CALC_SOFTMAX_LOOP_asn_1_itm_2;
      COMPUTE_BATCH_LOOP_asn_2_itm_3 <= COMPUTE_BATCH_LOOP_asn_2_itm_2;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_3 <= CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_2;
      CALC_SOFTMAX_LOOP_and_10_itm_3 <= CALC_SOFTMAX_LOOP_and_10_itm_2;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_3 <= exit_COMPUTE_BATCH_LOOP_sva_1_st_2;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_3 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( CALC_EXP_LOOP_and_6_cse ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_2 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_EXP_LOOP_and_svs_st_2 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_1_itm_2 <= 1'b0;
      COMPUTE_BATCH_LOOP_asn_2_itm_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_and_10_itm_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_2 <= 1'b0;
    end
    else if ( CALC_EXP_LOOP_and_6_cse ) begin
      CALC_EXP_LOOP_and_svs_st_2 <= CALC_EXP_LOOP_and_svs_st_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0;
      CALC_SOFTMAX_LOOP_asn_1_itm_2 <= CALC_SOFTMAX_LOOP_asn_1_itm_1;
      COMPUTE_BATCH_LOOP_asn_2_itm_2 <= exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_1;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_2 <= CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_1;
      CALC_SOFTMAX_LOOP_and_10_itm_2 <= CALC_SOFTMAX_LOOP_and_10_itm_1;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_2 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( CALC_SOFTMAX_LOOP_i_and_22_itm ) begin
      CALC_SOFTMAX_LOOP_i_7_0_lpi_1_6_0 <= MUX_v_7_2_2((signext_7_1(~ CALC_EXP_LOOP_and_svs_1)),
          (CALC_SOFTMAX_LOOP_acc_1_tmp[6:0]), CALC_SOFTMAX_LOOP_i_and_17_nl);
      SUM_EXP_LOOP_i_7_0_lpi_1_6_0 <= SUM_EXP_LOOP_acc_2_tmp[6:0];
      CALC_EXP_LOOP_i_7_0_lpi_1_6_0 <= CALC_EXP_LOOP_acc_1_tmp[6:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      COMPUTE_BATCH_LOOP_stage_0_7 <= 1'b0;
    end
    else if ( compute_wen & ((fsm_output[0]) | COMPUTE_BATCH_LOOP_stage_0_7_mx0c1)
        ) begin
      COMPUTE_BATCH_LOOP_stage_0_7 <= COMPUTE_BATCH_LOOP_stage_0_6 & COMPUTE_BATCH_LOOP_stage_0_7_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      COMPUTE_BATCH_LOOP_stage_0_8 <= 1'b0;
    end
    else if ( compute_wen & ((fsm_output[0]) | COMPUTE_BATCH_LOOP_stage_0_8_mx0c1)
        ) begin
      COMPUTE_BATCH_LOOP_stage_0_8 <= COMPUTE_BATCH_LOOP_stage_0_7 & COMPUTE_BATCH_LOOP_stage_0_8_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_COMPUTE_BATCH_LOOP_sva_1_st <= 1'b0;
    end
    else if ( compute_wen & CALC_SOFTMAX_LOOP_asn_itm & COMPUTE_BATCH_LOOP_and_33_tmp
        ) begin
      exit_COMPUTE_BATCH_LOOP_sva_1_st <= ~ COMPUTE_BATCH_LOOP_acc_itm_32_1;
    end
  end
  always @(posedge clk) begin
    if ( COMPUTE_BATCH_LOOP_and_64_cse ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_6 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_COMPUTE_BATCH_LOOP_sva_1_st_6 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_6 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_6 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_6 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0 <= 1'b0;
    end
    else if ( COMPUTE_BATCH_LOOP_and_64_cse ) begin
      exit_COMPUTE_BATCH_LOOP_sva_1_st_6 <= exit_COMPUTE_BATCH_LOOP_sva_1_st_5;
      CALC_SOFTMAX_LOOP_asn_itm_6 <= CALC_SOFTMAX_LOOP_asn_itm_5;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_6 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_5;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_6 <= exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_5;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_0;
    end
  end
  always @(posedge clk) begin
    if ( ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_and_cse
        ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm_1
          <= MUX_v_11_2_2(ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm_mx0w1,
          ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm,
          or_tmp_431);
      ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_9_0_itm_1
          <= MUX_v_10_2_2((ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[9:0]),
          ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_9_0_itm,
          or_tmp_431);
      ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm_1 <= MUX_v_8_2_2(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm_mx0w1,
          ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm, or_tmp_431);
    end
  end
  always @(posedge clk) begin
    if ( ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_and_cse ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_5 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_itm_1
          <= 1'b0;
      CALC_SOFTMAX_LOOP_and_10_itm_5 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_5 <= 1'b0;
    end
    else if ( ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_and_cse ) begin
      ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_itm_1
          <= ~((SUM_EXP_LOOP_acc_1_tmp!=74'b00000000000000000000000000000000000000000000000000000000000000000000000000));
      CALC_SOFTMAX_LOOP_and_10_itm_5 <= CALC_SOFTMAX_LOOP_and_10_itm_4;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_5 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( COMPUTE_BATCH_LOOP_and_65_cse ) begin
      CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_1 <= CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_2_6_0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_3 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_COMPUTE_BATCH_LOOP_sva_1_3 <= 1'b0;
    end
    else if ( COMPUTE_BATCH_LOOP_and_65_cse ) begin
      exit_COMPUTE_BATCH_LOOP_sva_1_3 <= exit_COMPUTE_BATCH_LOOP_sva_1_2;
    end
  end
  always @(posedge clk) begin
    if ( compute_wen & ((and_dcpl_165 & (fsm_output[1])) | CALC_EXP_LOOP_i_and_2_rgt)
        ) begin
      CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_1_6_0 <= MUX_v_7_2_2((signext_7_1(~ COMPUTE_BATCH_LOOP_acc_itm_32_1)),
          CALC_EXP_LOOP_i_7_0_lpi_1_6_0, CALC_EXP_LOOP_i_and_2_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_EXP_LOOP_and_svs_st_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_1_itm_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_and_10_itm_1 <= 1'b0;
    end
    else if ( CALC_EXP_LOOP_and_7_itm ) begin
      CALC_EXP_LOOP_and_svs_st_1 <= MUX_s_1_2_2(CALC_EXP_LOOP_and_svs_1, CALC_EXP_LOOP_and_svs_st,
          and_375_nl);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1, and_dcpl_166);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_0, and_dcpl_166);
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_1 <= (~ COMPUTE_BATCH_LOOP_acc_itm_32_1)
          & exitL_exit_CALC_SOFTMAX_LOOP_sva;
      CALC_SOFTMAX_LOOP_asn_1_itm_1 <= exitL_exit_CALC_SOFTMAX_LOOP_sva;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_or_tmp_1,
          CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm, and_dcpl_166);
      CALC_SOFTMAX_LOOP_and_10_itm_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_and_5_ssc_1,
          CALC_SOFTMAX_LOOP_and_10_itm, and_dcpl_166);
    end
  end
  always @(posedge clk) begin
    if ( ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_and_cse ) begin
      ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm <= ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm_mx0w1;
      ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_9_0_itm
          <= ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[9:0];
      ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm
          <= ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm_mx0w1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_COMPUTE_BATCH_LOOP_sva_1_2 <= 1'b0;
    end
    else if ( compute_wen & COMPUTE_BATCH_LOOP_and_28_tmp & (fsm_output[1]) ) begin
      exit_COMPUTE_BATCH_LOOP_sva_1_2 <= exit_COMPUTE_BATCH_LOOP_sva_1_1;
    end
  end
  always @(posedge clk) begin
    if ( compute_wen & CALC_EXP_LOOP_i_and_3_cse ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_2 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_EXP_LOOP_and_svs_st <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_31_cse & mux_141_cse & COMPUTE_BATCH_LOOP_and_33_tmp
        ) begin
      CALC_EXP_LOOP_and_svs_st <= CALC_EXP_LOOP_and_svs_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_0 <= 1'b0;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm <= 1'b0;
      CALC_SOFTMAX_LOOP_and_10_itm <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_89_cse ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm <= CALC_SOFTMAX_LOOP_or_tmp_1;
      CALC_SOFTMAX_LOOP_and_10_itm <= CALC_SOFTMAX_LOOP_and_5_ssc_1;
    end
  end
  always @(posedge clk) begin
    if ( COMPUTE_BATCH_LOOP_and_72_cse ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_1 <= CALC_SOFTMAX_LOOP_i_7_0_lpi_1_6_0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_COMPUTE_BATCH_LOOP_sva_1_1 <= 1'b0;
    end
    else if ( COMPUTE_BATCH_LOOP_and_72_cse ) begin
      exit_COMPUTE_BATCH_LOOP_sva_1_1 <= ~ COMPUTE_BATCH_LOOP_acc_itm_32_1;
    end
  end
  always @(posedge clk) begin
    if ( CALC_SOFTMAX_LOOP_i_and_34_cse ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_1 <= MUX_v_7_2_2(CALC_SOFTMAX_LOOP_i_7_0_lpi_1_6_0,
          CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm, and_dcpl_301);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_1 <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_i_and_34_cse ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_1 <= MUX_s_1_2_2((CALC_SOFTMAX_LOOP_acc_1_tmp[7]),
          CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm, and_dcpl_301);
    end
  end
  always @(posedge clk) begin
    if ( CALC_SOFTMAX_LOOP_i_and_36_cse ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm <= CALC_SOFTMAX_LOOP_i_7_0_lpi_1_6_0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_i_and_36_cse ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm <= CALC_SOFTMAX_LOOP_acc_1_tmp[7];
    end
  end
  assign nl_COMPUTE_BATCH_LOOP_acc_1_nl = COMPUTE_BATCH_LOOP_b_sva + 32'b00000000000000000000000000000001;
  assign COMPUTE_BATCH_LOOP_acc_1_nl = nl_COMPUTE_BATCH_LOOP_acc_1_nl[31:0];
  assign COMPUTE_BATCH_LOOP_b_and_nl = (or_dcpl_45 | (~ (CALC_SOFTMAX_LOOP_acc_1_tmp[7]))
      | exitL_exit_CALC_SOFTMAX_LOOP_sva | (~ COMPUTE_BATCH_LOOP_and_33_tmp)) & (fsm_output[1]);
  assign COMPUTE_BATCH_LOOP_b_mux_nl = MUX_v_32_2_2(COMPUTE_BATCH_LOOP_acc_1_nl,
      COMPUTE_BATCH_LOOP_b_sva, COMPUTE_BATCH_LOOP_b_and_nl);
  assign and_201_nl = nand_tmp_12 & COMPUTE_BATCH_LOOP_stage_0 & COMPUTE_BATCH_LOOP_and_33_tmp;
  assign and_203_nl = COMPUTE_BATCH_LOOP_stage_0 & (~ COMPUTE_BATCH_LOOP_stage_v);
  assign COMPUTE_BATCH_LOOP_mux1h_nl = MUX1HOT_s_1_3_2(exitL_exit_CALC_SOFTMAX_LOOP_sva_mx1w0,
      exitL_exit_CALC_SOFTMAX_LOOP_sva, CALC_SOFTMAX_LOOP_asn_itm, {and_201_nl ,
      and_203_nl , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_nand_1_cse});
  assign or_240_nl = and_dcpl_125 | (~ COMPUTE_BATCH_LOOP_and_33_tmp);
  assign COMPUTE_BATCH_LOOP_mux_86_nl = MUX_s_1_2_2(exitL_exit_CALC_SOFTMAX_LOOP_sva_mx1w0,
      exitL_exit_CALC_SOFTMAX_LOOP_sva, or_240_nl);
  assign and_nl = (~(or_cse & COMPUTE_BATCH_LOOP_stage_0_9)) & mux_21_cse;
  assign mux_292_nl = MUX_s_1_2_2(mux_21_cse, and_nl, or_8_cse);
  assign mux_293_nl = MUX_s_1_2_2(mux_21_cse, mux_292_nl, COMPUTE_BATCH_LOOP_stage_v_8);
  assign and_810_nl = nor_3_cse & (~(or_181_cse & plm_out_cnsi_bawt)) & or_120_cse;
  assign mux_302_nl = MUX_s_1_2_2(or_120_cse, and_810_nl, and_dcpl_147);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_2_nl
      = MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28[11:10]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_3_nl
      = MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28[11:10]);
  assign nl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:10])
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_2_nl
      , 1'b1 , ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_3_nl});
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign operator_74_54_false_AC_TRN_AC_WRAP_1_mux_nl = MUX_s_1_2_2(COMPUTE_BATCH_LOOP_stage_0_1,
      COMPUTE_BATCH_LOOP_stage_0, COMPUTE_BATCH_LOOP_and_33_tmp);
  assign nor_125_nl = ~(COMPUTE_BATCH_LOOP_and_28_tmp | COMPUTE_BATCH_LOOP_and_33_tmp);
  assign COMPUTE_BATCH_LOOP_mux_85_nl = MUX_s_1_2_2(COMPUTE_BATCH_LOOP_stage_0_1,
      COMPUTE_BATCH_LOOP_stage_0_2, nor_125_nl);
  assign nor_126_nl = ~(COMPUTE_BATCH_LOOP_and_23_tmp | COMPUTE_BATCH_LOOP_and_28_tmp);
  assign COMPUTE_BATCH_LOOP_mux_84_nl = MUX_s_1_2_2(COMPUTE_BATCH_LOOP_stage_0_2,
      COMPUTE_BATCH_LOOP_stage_0_3, nor_126_nl);
  assign nor_122_nl = ~(COMPUTE_BATCH_LOOP_and_23_tmp | COMPUTE_BATCH_LOOP_and_19_tmp);
  assign COMPUTE_BATCH_LOOP_mux_83_nl = MUX_s_1_2_2(COMPUTE_BATCH_LOOP_stage_0_3,
      COMPUTE_BATCH_LOOP_stage_0_4, nor_122_nl);
  assign nor_123_nl = ~(COMPUTE_BATCH_LOOP_and_19_tmp | COMPUTE_BATCH_LOOP_and_16_tmp);
  assign COMPUTE_BATCH_LOOP_mux_82_nl = MUX_s_1_2_2(COMPUTE_BATCH_LOOP_stage_0_4,
      COMPUTE_BATCH_LOOP_stage_0_5, nor_123_nl);
  assign nor_124_nl = ~(COMPUTE_BATCH_LOOP_and_16_tmp | COMPUTE_BATCH_LOOP_and_13_tmp);
  assign COMPUTE_BATCH_LOOP_mux_81_nl = MUX_s_1_2_2(COMPUTE_BATCH_LOOP_stage_0_5,
      COMPUTE_BATCH_LOOP_stage_0_6, nor_124_nl);
  assign nor_94_nl = ~(COMPUTE_BATCH_LOOP_stage_v_8 | (~ and_tmp_85));
  assign mux_281_nl = MUX_s_1_2_2(and_tmp_85, and_244_cse, COMPUTE_BATCH_LOOP_stage_v_8);
  assign mux_282_nl = MUX_s_1_2_2(nor_94_nl, mux_281_nl, or_8_cse);
  assign COMPUTE_BATCH_LOOP_mux_80_nl = MUX_s_1_2_2(COMPUTE_BATCH_LOOP_stage_0_9,
      COMPUTE_BATCH_LOOP_stage_0_8, mux_282_nl);
  assign and_264_nl = or_48_cse & COMPUTE_BATCH_LOOP_stage_v_8 & COMPUTE_BATCH_LOOP_stage_0_9
      & or_106_cse;
  assign and_263_nl = or_46_cse & COMPUTE_BATCH_LOOP_stage_v_8 & COMPUTE_BATCH_LOOP_stage_0_9
      & or_106_cse;
  assign mux_295_nl = MUX_s_1_2_2(and_264_nl, and_263_nl, plm_out_cnsi_bawt);
  assign nand_20_nl = ~(or_cse & or_8_cse & mux_295_nl);
  assign nand_21_nl = ~(COMPUTE_BATCH_LOOP_stage_0_10 & mux_271_cse);
  assign mux_296_nl = MUX_s_1_2_2(nand_20_nl, nand_21_nl, reg_COMPUTE_BATCH_LOOP_stage_v_9_cse);
  assign COMPUTE_BATCH_LOOP_mux_79_nl = MUX_s_1_2_2(COMPUTE_BATCH_LOOP_stage_0_9,
      COMPUTE_BATCH_LOOP_stage_0_10, mux_296_nl);
  assign and_284_nl = CALC_SOFTMAX_LOOP_asn_itm & COMPUTE_BATCH_LOOP_and_33_tmp;
  assign and_285_nl = (~ CALC_SOFTMAX_LOOP_asn_itm) & COMPUTE_BATCH_LOOP_and_33_tmp;
  assign CALC_SOFTMAX_LOOP_i_and_17_nl = CALC_SOFTMAX_LOOP_equal_tmp_2 & COMPUTE_BATCH_LOOP_and_33_tmp;
  assign and_375_nl = (~ mux_141_cse) & COMPUTE_BATCH_LOOP_and_33_tmp;

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [73:0] MUX1HOT_v_74_3_2;
    input [73:0] input_2;
    input [73:0] input_1;
    input [73:0] input_0;
    input [2:0] sel;
    reg [73:0] result;
  begin
    result = input_0 & {74{sel[0]}};
    result = result | ( input_1 & {74{sel[1]}});
    result = result | ( input_2 & {74{sel[2]}});
    MUX1HOT_v_74_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_8_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [9:0] input_2;
    input [9:0] input_3;
    input [9:0] input_4;
    input [9:0] input_5;
    input [9:0] input_6;
    input [9:0] input_7;
    input [2:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_10_8_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_4_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [1:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_3_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_4_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [4:0] input_2;
    input [4:0] input_3;
    input [1:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_5_4_2 = result;
  end
  endfunction


  function automatic [66:0] MUX_v_67_2_2;
    input [66:0] input_0;
    input [66:0] input_1;
    input [0:0] sel;
    reg [66:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_67_2_2 = result;
  end
  endfunction


  function automatic [73:0] MUX_v_74_2_2;
    input [73:0] input_0;
    input [73:0] input_1;
    input [0:0] sel;
    reg [73:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_74_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_4_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [6:0] input_2;
    input [6:0] input_3;
    input [1:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_7_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_8_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2 = result;
  end
  endfunction


  function automatic [93:0] MUX_v_94_2_2;
    input [93:0] input_0;
    input [93:0] input_1;
    input [0:0] sel;
    reg [93:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_94_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [18:0] readslicef_47_19_28;
    input [46:0] vector;
    reg [46:0] tmp;
  begin
    tmp = vector >> 28;
    readslicef_47_19_28 = tmp[18:0];
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input [0:0] vector;
  begin
    signext_7_1= {{6{vector[0]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_s2u_9_11 = {{2{vector[8]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_11 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [18:0] conv_u2u_19_19 ;
    input [18:0]  vector ;
  begin
    conv_u2u_19_19 = vector;
  end
  endfunction


  function automatic [32:0] conv_u2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_33 = {1'b0, vector};
  end
  endfunction


  function automatic [73:0] conv_u2u_67_74 ;
    input [66:0]  vector ;
  begin
    conv_u2u_67_74 = {{7{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load_load
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load_load (
  clk, rst, conf_info, dma_read_ctrl_val, dma_read_ctrl_rdy, dma_read_ctrl_msg, dma_read_chnl_val,
      dma_read_chnl_rdy, dma_read_chnl_msg, done, input_ready_req_req, input_ready_ack_ack,
      plm_in_cns_req_vz, plm_in_cns_rls_lz, plm_in_cnsi_d_d, plm_in_cnsi_wadr_d,
      plm_in_cnsi_we_d_pff
);
  input clk;
  input rst;
  input [31:0] conf_info;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  input done;
  output input_ready_req_req;
  input input_ready_ack_ack;
  input plm_in_cns_req_vz;
  output plm_in_cns_rls_lz;
  output [31:0] plm_in_cnsi_d_d;
  output [6:0] plm_in_cnsi_wadr_d;
  output plm_in_cnsi_we_d_pff;


  // Interconnect Declarations
  wire load_wen;
  wire dma_read_ctrl_Push_mioi_bawt;
  reg dma_read_ctrl_Push_mioi_iswt0;
  wire load_wten;
  wire dma_read_ctrl_Push_mioi_wen_comp;
  reg dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_psct;
  wire dma_read_chnl_Pop_mioi_bawt;
  reg dma_read_chnl_Pop_mioi_iswt0;
  wire dma_read_chnl_Pop_mioi_wen_comp;
  wire [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt;
  reg dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_psct;
  wire input_ready_req_mioi_bawt;
  wire input_ready_req_mioi_wen_comp;
  reg input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_psct;
  wire plm_in_cnsi_bawt;
  wire plm_in_cns_rls_obj_bawt;
  wire plm_in_cns_req_obj_bawt;
  reg plm_in_cns_req_obj_iswt0;
  wire plm_in_cns_req_obj_wen_comp;
  reg [3:0] dma_read_ctrl_Push_mioi_m_index_rsc_dat_10_7;
  wire [2:0] fsm_output;
  wire [4:0] LOAD_BATCH_LOOP_acc_2_tmp;
  wire [5:0] nl_LOAD_BATCH_LOOP_acc_2_tmp;
  wire [7:0] LOAD_LOOP_acc_2_tmp;
  wire [8:0] nl_LOAD_LOOP_acc_2_tmp;
  wire LOAD_BATCH_LOOP_and_8_tmp;
  wire LOAD_BATCH_LOOP_and_4_tmp;
  wire or_dcpl_5;
  wire and_dcpl_4;
  wire and_dcpl_6;
  wire or_dcpl_18;
  wire and_dcpl_11;
  wire and_dcpl_14;
  wire and_dcpl_15;
  wire and_dcpl_17;
  wire or_dcpl_22;
  wire or_dcpl_23;
  wire and_dcpl_25;
  wire or_dcpl_27;
  wire or_dcpl_30;
  wire or_tmp_35;
  wire mux_tmp_41;
  wire mux_tmp_42;
  wire or_dcpl_41;
  wire and_dcpl_56;
  wire or_tmp_38;
  wire or_tmp_39;
  wire or_tmp_44;
  wire or_tmp_46;
  wire or_tmp_59;
  reg exitL_exit_LOAD_LOOP_sva;
  reg LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_2;
  reg LOAD_BATCH_LOOP_stage_v_2;
  reg LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_3;
  reg exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_3;
  reg LOAD_BATCH_LOOP_stage_v_3;
  reg exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_1;
  reg LOAD_BATCH_LOOP_stage_0_3;
  reg LOAD_LOOP_asn_itm;
  reg LOAD_BATCH_LOOP_stage_0;
  reg exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2;
  reg LOAD_BATCH_LOOP_stage_0_1;
  reg LOAD_BATCH_LOOP_stage_0_2;
  reg LOAD_BATCH_LOOP_stage_v;
  reg exit_LOAD_BATCH_LOOP_sva_1_st_1;
  reg LOAD_LOOP_asn_itm_1;
  reg LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_1;
  reg reg_dma_read_chnl_Pop_mioi_oswt_cse;
  reg reg_input_ready_req_mioi_iswt0_cse;
  reg reg_plm_in_cns_rls_obj_iswt0_cse;
  wire and_162_cse;
  wire LOAD_LOOP_i_and_cse;
  wire LOAD_LOOP_LOAD_LOOP_and_cse;
  wire or_57_cse;
  reg [31:0] plm_in_cnsi_d_d_reg;
  wire [31:0] LOAD_LOOP_mux_rmff;
  reg [6:0] plm_in_cnsi_wadr_d_reg;
  wire [6:0] LOAD_LOOP_i_mux_rmff;
  wire plm_in_cnsi_we_d_iff;
  wire and_74_rmff;
  wire and_70_rmff;
  wire [3:0] LOAD_BATCH_LOOP_b_mux_rmff;
  wire LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_or_2_rmff;
  wire LOAD_LOOP_LOAD_LOOP_or_rmff;
  wire softmax_sysc_load_compute_handshake_softmax_sysc_load_compute_handshake_or_rmff;
  wire LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_and_itm;
  reg [31:0] config_batch_sva;
  reg LOAD_BATCH_LOOP_stage_v_1;
  reg exit_LOAD_BATCH_LOOP_sva_1_st;
  reg LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm;
  reg [6:0] LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_6_0_itm_1;
  reg [6:0] LOAD_LOOP_i_7_0_lpi_1_6_0;
  reg [3:0] LOAD_BATCH_LOOP_b_4_0_sva_3_0;
  wire exitL_exit_LOAD_LOOP_sva_mx1w0;
  wire LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_or_cse_1;
  wire LOAD_BATCH_LOOP_nand_12_cse_1;
  wire and_60_rgt;
  wire LOAD_BATCH_LOOP_acc_1_itm_32_1;

  wire[0:0] or_99_nl;
  wire[3:0] LOAD_BATCH_LOOP_b_mux_2_nl;
  wire[0:0] LOAD_BATCH_LOOP_b_and_nl;
  wire[0:0] LOAD_BATCH_LOOP_mux1h_nl;
  wire[0:0] and_42_nl;
  wire[0:0] and_44_nl;
  wire[0:0] or_74_nl;
  wire[0:0] LOAD_BATCH_LOOP_mux_26_nl;
  wire[0:0] or_76_nl;
  wire[0:0] and_57_nl;
  wire[0:0] and_58_nl;
  wire[0:0] LOAD_LOOP_i_nand_nl;
  wire[0:0] LOAD_LOOP_i_and_4_nl;
  wire[0:0] and_61_nl;
  wire[0:0] LOAD_BATCH_LOOP_mux_23_nl;
  wire[0:0] LOAD_BATCH_LOOP_mux_25_nl;
  wire[0:0] nor_nl;
  wire[0:0] LOAD_BATCH_LOOP_mux_24_nl;
  wire[0:0] and_48_nl;
  wire[32:0] LOAD_BATCH_LOOP_acc_1_nl;
  wire[33:0] nl_LOAD_BATCH_LOOP_acc_1_nl;
  wire[6:0] LOAD_LOOP_mux_5_nl;
  wire[0:0] and_45_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_softmax_sysc_load_load_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat;
  assign nl_softmax_sysc_load_load_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat
      = {21'b000000000000000000000 , LOAD_BATCH_LOOP_b_mux_rmff , 7'b0000000};
  wire [0:0] nl_softmax_sysc_load_load_input_ready_req_mioi_inst_input_ready_req_mioi_oswt_unreg;
  assign nl_softmax_sysc_load_load_input_ready_req_mioi_inst_input_ready_req_mioi_oswt_unreg
      = and_dcpl_17 & (fsm_output[1]);
  wire [0:0] nl_softmax_sysc_load_load_plm_in_cnsi_1_inst_plm_in_cnsi_oswt_unreg;
  assign nl_softmax_sysc_load_load_plm_in_cnsi_1_inst_plm_in_cnsi_oswt_unreg = or_dcpl_23
      & or_57_cse & and_dcpl_25 & plm_in_cnsi_bawt & (~ exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2)
      & (fsm_output[1]);
  wire [0:0] nl_softmax_sysc_load_load_load_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  assign nl_softmax_sysc_load_load_load_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0 = ~
      done;
  wire [0:0] nl_softmax_sysc_load_load_load_fsm_inst_LOAD_BATCH_LOOP_C_0_tr0;
  assign nl_softmax_sysc_load_load_load_fsm_inst_LOAD_BATCH_LOOP_C_0_tr0 = LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_and_itm
      | (~((~(and_dcpl_4 & (~ input_ready_req_mioi_bawt))) & LOAD_BATCH_LOOP_stage_v_3))
      | LOAD_BATCH_LOOP_stage_0_3 | LOAD_BATCH_LOOP_stage_0_2 | LOAD_BATCH_LOOP_stage_0_1;
  esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_ctrl_Push_mioi softmax_sysc_load_load_dma_read_ctrl_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_ctrl_val(dma_read_ctrl_val),
      .dma_read_ctrl_rdy(dma_read_ctrl_rdy),
      .dma_read_ctrl_msg(dma_read_ctrl_msg),
      .load_wen(load_wen),
      .dma_read_ctrl_Push_mioi_m_index_rsc_dat(nl_softmax_sysc_load_load_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat[31:0]),
      .dma_read_ctrl_Push_mioi_oswt_unreg(and_70_rmff),
      .dma_read_ctrl_Push_mioi_bawt(dma_read_ctrl_Push_mioi_bawt),
      .dma_read_ctrl_Push_mioi_iswt0(dma_read_ctrl_Push_mioi_iswt0),
      .load_wten(load_wten),
      .dma_read_ctrl_Push_mioi_wen_comp(dma_read_ctrl_Push_mioi_wen_comp),
      .dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_psct(LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_or_2_rmff),
      .dma_read_ctrl_Push_mioi_iswt0_pff(or_tmp_38)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_dma_read_chnl_Pop_mioi softmax_sysc_load_load_dma_read_chnl_Pop_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_chnl_val(dma_read_chnl_val),
      .dma_read_chnl_rdy(dma_read_chnl_rdy),
      .dma_read_chnl_msg(dma_read_chnl_msg),
      .load_wen(load_wen),
      .load_wten(load_wten),
      .dma_read_chnl_Pop_mioi_oswt_unreg(and_74_rmff),
      .dma_read_chnl_Pop_mioi_bawt(dma_read_chnl_Pop_mioi_bawt),
      .dma_read_chnl_Pop_mioi_iswt0(dma_read_chnl_Pop_mioi_iswt0),
      .dma_read_chnl_Pop_mioi_wen_comp(dma_read_chnl_Pop_mioi_wen_comp),
      .dma_read_chnl_Pop_mioi_return_rsc_z_mxwt(dma_read_chnl_Pop_mioi_return_rsc_z_mxwt),
      .dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_psct(LOAD_LOOP_LOAD_LOOP_or_rmff),
      .dma_read_chnl_Pop_mioi_iswt0_pff(or_tmp_44)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_input_ready_req_mioi softmax_sysc_load_load_input_ready_req_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .input_ready_req_req(input_ready_req_req),
      .input_ready_ack_ack(input_ready_ack_ack),
      .load_wen(load_wen),
      .load_wten(load_wten),
      .input_ready_req_mioi_oswt_unreg(nl_softmax_sysc_load_load_input_ready_req_mioi_inst_input_ready_req_mioi_oswt_unreg[0:0]),
      .input_ready_req_mioi_bawt(input_ready_req_mioi_bawt),
      .input_ready_req_mioi_iswt0(reg_input_ready_req_mioi_iswt0_cse),
      .input_ready_req_mioi_wen_comp(input_ready_req_mioi_wen_comp),
      .input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_psct(softmax_sysc_load_compute_handshake_softmax_sysc_load_compute_handshake_or_rmff),
      .input_ready_req_mioi_iswt0_pff(or_tmp_46)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cnsi_1 softmax_sysc_load_load_plm_in_cnsi_1_inst
      (
      .clk(clk),
      .rst(rst),
      .load_wen(load_wen),
      .load_wten(load_wten),
      .plm_in_cnsi_oswt_unreg(nl_softmax_sysc_load_load_plm_in_cnsi_1_inst_plm_in_cnsi_oswt_unreg[0:0]),
      .plm_in_cnsi_bawt(plm_in_cnsi_bawt),
      .plm_in_cnsi_iswt0(reg_dma_read_chnl_Pop_mioi_oswt_cse),
      .plm_in_cnsi_we_d_pff(plm_in_cnsi_we_d_iff),
      .plm_in_cnsi_iswt0_pff(and_74_rmff)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_rls_obj softmax_sysc_load_load_plm_in_cns_rls_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_rls_lz(plm_in_cns_rls_lz),
      .load_wen(load_wen),
      .load_wten(load_wten),
      .plm_in_cns_rls_obj_oswt_unreg(or_tmp_46),
      .plm_in_cns_rls_obj_bawt(plm_in_cns_rls_obj_bawt),
      .plm_in_cns_rls_obj_iswt0(reg_plm_in_cns_rls_obj_iswt0_cse)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_plm_in_cns_req_obj softmax_sysc_load_load_plm_in_cns_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_req_vz(plm_in_cns_req_vz),
      .load_wen(load_wen),
      .plm_in_cns_req_obj_oswt_unreg(and_70_rmff),
      .plm_in_cns_req_obj_bawt(plm_in_cns_req_obj_bawt),
      .plm_in_cns_req_obj_iswt0(plm_in_cns_req_obj_iswt0),
      .plm_in_cns_req_obj_wen_comp(plm_in_cns_req_obj_wen_comp)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_staller softmax_sysc_load_load_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .load_wen(load_wen),
      .load_wten(load_wten),
      .dma_read_ctrl_Push_mioi_wen_comp(dma_read_ctrl_Push_mioi_wen_comp),
      .dma_read_chnl_Pop_mioi_wen_comp(dma_read_chnl_Pop_mioi_wen_comp),
      .input_ready_req_mioi_wen_comp(input_ready_req_mioi_wen_comp),
      .plm_in_cns_req_obj_wen_comp(plm_in_cns_req_obj_wen_comp)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load_load_fsm softmax_sysc_load_load_load_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .load_wen(load_wen),
      .fsm_output(fsm_output),
      .WAIT_FOR_CONFIG_LOOP_C_0_tr0(nl_softmax_sysc_load_load_load_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0[0:0]),
      .LOAD_BATCH_LOOP_C_0_tr0(nl_softmax_sysc_load_load_load_fsm_inst_LOAD_BATCH_LOOP_C_0_tr0[0:0])
    );
  assign and_70_rmff = and_dcpl_11 & (fsm_output[1]);
  assign and_74_rmff = and_dcpl_14 & (fsm_output[1]);
  assign or_57_cse = plm_in_cns_rls_obj_bawt | (~ LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_2);
  assign softmax_sysc_load_compute_handshake_softmax_sysc_load_compute_handshake_or_rmff
      = (input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_psct & (~((or_dcpl_27
      | (~ plm_in_cnsi_bawt) | (~ plm_in_cns_rls_obj_bawt) | (~ LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_2)
      | exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2) & and_dcpl_17 & (fsm_output[1])))) |
      or_tmp_46;
  assign or_99_nl = or_dcpl_18 | (~ (fsm_output[1]));
  assign LOAD_BATCH_LOOP_b_mux_rmff = MUX_v_4_2_2(LOAD_BATCH_LOOP_b_4_0_sva_3_0,
      dma_read_ctrl_Push_mioi_m_index_rsc_dat_10_7, or_99_nl);
  assign LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_or_2_rmff = (dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_psct
      & (~ or_tmp_39)) | or_tmp_38;
  assign LOAD_LOOP_LOAD_LOOP_or_rmff = (dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_psct
      & (~(or_dcpl_30 & and_dcpl_14 & (fsm_output[1])))) | or_tmp_44;
  assign LOAD_LOOP_i_mux_rmff = MUX_v_7_2_2(LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_6_0_itm_1,
      plm_in_cnsi_wadr_d_reg, or_tmp_59);
  assign LOAD_LOOP_mux_rmff = MUX_v_32_2_2(dma_read_chnl_Pop_mioi_return_rsc_z_mxwt,
      plm_in_cnsi_d_d_reg, or_tmp_59);
  assign LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_and_itm = LOAD_BATCH_LOOP_stage_0 & (and_dcpl_6
      | (~ LOAD_BATCH_LOOP_and_8_tmp));
  assign and_162_cse = (LOAD_LOOP_acc_2_tmp[7]) & (LOAD_BATCH_LOOP_acc_2_tmp[4]);
  assign LOAD_LOOP_i_and_cse = load_wen & (fsm_output[1]);
  assign and_60_rgt = (~ LOAD_BATCH_LOOP_acc_1_itm_32_1) & and_dcpl_56;
  assign LOAD_LOOP_LOAD_LOOP_and_cse = (~ LOAD_BATCH_LOOP_acc_1_itm_32_1) & exitL_exit_LOAD_LOOP_sva;
  assign exitL_exit_LOAD_LOOP_sva_mx1w0 = ~((LOAD_BATCH_LOOP_acc_2_tmp[4]) | (~ (LOAD_LOOP_acc_2_tmp[7])));
  assign nl_LOAD_BATCH_LOOP_acc_1_nl = ({29'b10000000000000000000000000000 , LOAD_BATCH_LOOP_b_4_0_sva_3_0})
      + conv_u2u_32_33(~ config_batch_sva) + 33'b000000000000000000000000000000001;
  assign LOAD_BATCH_LOOP_acc_1_nl = nl_LOAD_BATCH_LOOP_acc_1_nl[32:0];
  assign LOAD_BATCH_LOOP_acc_1_itm_32_1 = readslicef_33_1_32(LOAD_BATCH_LOOP_acc_1_nl);
  assign nl_LOAD_BATCH_LOOP_acc_2_tmp = conv_u2u_4_5(LOAD_BATCH_LOOP_b_4_0_sva_3_0)
      + 5'b00001;
  assign LOAD_BATCH_LOOP_acc_2_tmp = nl_LOAD_BATCH_LOOP_acc_2_tmp[4:0];
  assign LOAD_LOOP_mux_5_nl = MUX_v_7_2_2(LOAD_LOOP_i_7_0_lpi_1_6_0, (signext_7_1(~
      LOAD_BATCH_LOOP_acc_1_itm_32_1)), exitL_exit_LOAD_LOOP_sva);
  assign nl_LOAD_LOOP_acc_2_tmp = conv_u2u_7_8(LOAD_LOOP_mux_5_nl) + 8'b00000001;
  assign LOAD_LOOP_acc_2_tmp = nl_LOAD_LOOP_acc_2_tmp[7:0];
  assign LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_or_cse_1 = input_ready_req_mioi_bawt | (~(LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_3
      & (~ exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_3) & LOAD_BATCH_LOOP_stage_v_3));
  assign LOAD_BATCH_LOOP_nand_12_cse_1 = ~((~ exit_LOAD_BATCH_LOOP_sva_1_st_1) &
      LOAD_LOOP_asn_itm_1 & LOAD_BATCH_LOOP_stage_v_1);
  assign LOAD_BATCH_LOOP_and_8_tmp = LOAD_BATCH_LOOP_stage_v & (~(LOAD_BATCH_LOOP_stage_v_1
      & (~ LOAD_BATCH_LOOP_and_4_tmp))) & LOAD_BATCH_LOOP_stage_0_1 & (plm_in_cnsi_bawt
      | (~((~ exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2) & LOAD_BATCH_LOOP_stage_v_2)))
      & (plm_in_cns_rls_obj_bawt | (~(LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_2 & (~
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2) & LOAD_BATCH_LOOP_stage_v_2))) & LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_or_cse_1;
  assign LOAD_BATCH_LOOP_and_4_tmp = LOAD_BATCH_LOOP_stage_v_1 & (~(LOAD_BATCH_LOOP_stage_v_2
      & or_dcpl_41)) & LOAD_BATCH_LOOP_stage_0_2 & (dma_read_ctrl_Push_mioi_bawt
      | LOAD_BATCH_LOOP_nand_12_cse_1) & (plm_in_cns_req_obj_bawt | LOAD_BATCH_LOOP_nand_12_cse_1)
      & (dma_read_chnl_Pop_mioi_bawt | exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_1) & LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_or_cse_1;
  assign or_dcpl_5 = LOAD_BATCH_LOOP_acc_1_itm_32_1 | (~ exitL_exit_LOAD_LOOP_sva);
  assign and_dcpl_4 = LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_3 & (~ exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_3);
  assign and_dcpl_6 = or_dcpl_5 & (~((LOAD_BATCH_LOOP_acc_2_tmp[4]) & (LOAD_LOOP_acc_2_tmp[7])));
  assign or_dcpl_18 = ~(LOAD_BATCH_LOOP_acc_1_itm_32_1 & LOAD_LOOP_asn_itm & LOAD_BATCH_LOOP_and_8_tmp);
  assign and_dcpl_11 = LOAD_BATCH_LOOP_and_4_tmp & (~ exit_LOAD_BATCH_LOOP_sva_1_st_1)
      & LOAD_LOOP_asn_itm_1;
  assign and_dcpl_14 = LOAD_BATCH_LOOP_and_4_tmp & (~ exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_1);
  assign and_dcpl_15 = or_dcpl_5 & LOAD_BATCH_LOOP_and_8_tmp;
  assign and_dcpl_17 = and_dcpl_4 & input_ready_req_mioi_bawt & LOAD_BATCH_LOOP_stage_v_3;
  assign or_dcpl_22 = (~ LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_3) | exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_3;
  assign or_dcpl_23 = or_dcpl_22 | input_ready_req_mioi_bawt | (~ LOAD_BATCH_LOOP_stage_v_3);
  assign and_dcpl_25 = LOAD_BATCH_LOOP_stage_0_3 & LOAD_BATCH_LOOP_stage_v_2;
  assign or_dcpl_27 = ~(LOAD_BATCH_LOOP_stage_0_3 & LOAD_BATCH_LOOP_stage_v_2);
  assign or_dcpl_30 = LOAD_LOOP_LOAD_LOOP_and_cse | (~ LOAD_BATCH_LOOP_and_8_tmp);
  assign or_tmp_35 = and_162_cse | LOAD_LOOP_LOAD_LOOP_and_cse;
  assign mux_tmp_41 = MUX_s_1_2_2(LOAD_BATCH_LOOP_stage_v, or_tmp_35, LOAD_BATCH_LOOP_and_8_tmp);
  assign and_45_nl = or_57_cse & plm_in_cnsi_bawt & or_dcpl_23;
  assign mux_tmp_42 = MUX_s_1_2_2(and_45_nl, or_dcpl_23, exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2);
  assign or_dcpl_41 = (~ mux_tmp_42) | or_dcpl_27;
  assign and_dcpl_56 = exitL_exit_LOAD_LOOP_sva & LOAD_BATCH_LOOP_and_8_tmp;
  assign or_tmp_38 = LOAD_BATCH_LOOP_acc_1_itm_32_1 & LOAD_LOOP_asn_itm & LOAD_BATCH_LOOP_and_8_tmp
      & (fsm_output[1]);
  assign or_tmp_39 = and_dcpl_11 & or_dcpl_18 & (fsm_output[1]);
  assign or_tmp_44 = and_dcpl_15 & (fsm_output[1]);
  assign or_tmp_46 = or_dcpl_23 & LOAD_BATCH_LOOP_stage_0_3 & LOAD_BATCH_LOOP_stage_v_2
      & plm_in_cnsi_bawt & plm_in_cns_rls_obj_bawt & LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_2
      & (~ exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2) & (fsm_output[1]);
  assign or_tmp_59 = (~ LOAD_BATCH_LOOP_and_4_tmp) | exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_1
      | (~ (fsm_output[1]));
  assign plm_in_cnsi_d_d = LOAD_LOOP_mux_rmff;
  assign plm_in_cnsi_wadr_d = LOAD_LOOP_i_mux_rmff;
  assign plm_in_cnsi_we_d_pff = plm_in_cnsi_we_d_iff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cns_req_obj_iswt0 <= 1'b0;
    end
    else if ( load_wen & (or_tmp_38 | or_tmp_39) ) begin
      plm_in_cns_req_obj_iswt0 <= ~ or_tmp_39;
    end
  end
  always @(posedge clk) begin
    if ( load_wen ) begin
      input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_psct <= softmax_sysc_load_compute_handshake_softmax_sysc_load_compute_handshake_or_rmff;
      dma_read_ctrl_Push_mioi_m_index_rsc_dat_10_7 <= LOAD_BATCH_LOOP_b_mux_rmff;
      dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_psct <= LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_or_2_rmff;
      dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_psct <= LOAD_LOOP_LOAD_LOOP_or_rmff;
      plm_in_cnsi_wadr_d_reg <= LOAD_LOOP_i_mux_rmff;
      plm_in_cnsi_d_d_reg <= LOAD_LOOP_mux_rmff;
      LOAD_BATCH_LOOP_b_4_0_sva_3_0 <= MUX_v_4_2_2(4'b0000, LOAD_BATCH_LOOP_b_mux_2_nl,
          (fsm_output[1]));
      config_batch_sva <= MUX_v_32_2_2(conf_info, config_batch_sva, fsm_output[1]);
      LOAD_BATCH_LOOP_stage_v_1 <= ((LOAD_BATCH_LOOP_stage_v_1 & (~ LOAD_BATCH_LOOP_and_4_tmp))
          | LOAD_BATCH_LOOP_and_8_tmp) & (fsm_output[1]);
      LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_6_0_itm_1 <= MUX1HOT_v_7_3_2(LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_6_0_itm_1,
          (signext_7_1(~ LOAD_BATCH_LOOP_acc_1_itm_32_1)), LOAD_LOOP_i_7_0_lpi_1_6_0,
          {LOAD_LOOP_i_nand_nl , LOAD_LOOP_i_and_4_nl , and_61_nl});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_Push_mioi_iswt0 <= 1'b0;
      reg_dma_read_chnl_Pop_mioi_oswt_cse <= 1'b0;
      dma_read_chnl_Pop_mioi_iswt0 <= 1'b0;
      reg_input_ready_req_mioi_iswt0_cse <= 1'b0;
      reg_plm_in_cns_rls_obj_iswt0_cse <= 1'b0;
      LOAD_BATCH_LOOP_stage_v <= 1'b0;
      LOAD_BATCH_LOOP_stage_0 <= 1'b0;
      LOAD_LOOP_asn_itm <= 1'b0;
      exitL_exit_LOAD_LOOP_sva <= 1'b0;
      LOAD_BATCH_LOOP_stage_v_2 <= 1'b0;
      LOAD_BATCH_LOOP_stage_v_3 <= 1'b0;
      LOAD_BATCH_LOOP_stage_0_1 <= 1'b0;
      LOAD_BATCH_LOOP_stage_0_2 <= 1'b0;
      LOAD_BATCH_LOOP_stage_0_3 <= 1'b0;
    end
    else if ( load_wen ) begin
      dma_read_ctrl_Push_mioi_iswt0 <= or_tmp_38;
      reg_dma_read_chnl_Pop_mioi_oswt_cse <= and_74_rmff;
      dma_read_chnl_Pop_mioi_iswt0 <= or_tmp_44;
      reg_input_ready_req_mioi_iswt0_cse <= or_tmp_46;
      reg_plm_in_cns_rls_obj_iswt0_cse <= and_dcpl_14 & LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_1
          & (fsm_output[1]);
      LOAD_BATCH_LOOP_stage_v <= ~((~(LOAD_BATCH_LOOP_stage_v & (~((LOAD_LOOP_LOAD_LOOP_and_cse
          | and_162_cse | (~ LOAD_BATCH_LOOP_stage_0)) & LOAD_BATCH_LOOP_and_8_tmp))))
          & (~((~ mux_tmp_41) & LOAD_BATCH_LOOP_stage_0)) & (fsm_output[1]));
      LOAD_BATCH_LOOP_stage_0 <= LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_and_itm | (~ (fsm_output[1]));
      LOAD_LOOP_asn_itm <= LOAD_BATCH_LOOP_mux1h_nl | (~ (fsm_output[1]));
      exitL_exit_LOAD_LOOP_sva <= LOAD_BATCH_LOOP_mux_26_nl | (~ (fsm_output[1]));
      LOAD_BATCH_LOOP_stage_v_2 <= ((LOAD_BATCH_LOOP_stage_v_2 & (~(mux_tmp_42 &
          and_dcpl_25))) | LOAD_BATCH_LOOP_and_4_tmp) & (fsm_output[1]);
      LOAD_BATCH_LOOP_stage_v_3 <= ((LOAD_BATCH_LOOP_stage_v_3 & (~(((~(((~((~ plm_in_cns_rls_obj_bawt)
          & LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_2)) & plm_in_cnsi_bawt) | exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2))
          | or_dcpl_27) & (or_dcpl_22 | input_ready_req_mioi_bawt)))) | (mux_tmp_42
          & and_dcpl_25)) & (fsm_output[1]);
      LOAD_BATCH_LOOP_stage_0_1 <= ~((~(LOAD_BATCH_LOOP_mux_23_nl & (~(or_tmp_35
          & LOAD_BATCH_LOOP_and_8_tmp)))) & (fsm_output[1]));
      LOAD_BATCH_LOOP_stage_0_2 <= LOAD_BATCH_LOOP_mux_25_nl & (fsm_output[1]);
      LOAD_BATCH_LOOP_stage_0_3 <= LOAD_BATCH_LOOP_mux_24_nl & (fsm_output[1]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_2 <= 1'b0;
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2 <= 1'b0;
      LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_3 <= 1'b0;
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_3 <= 1'b0;
      exit_LOAD_BATCH_LOOP_sva_1_st_1 <= 1'b0;
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_1 <= 1'b0;
      LOAD_LOOP_asn_itm_1 <= 1'b0;
    end
    else if ( LOAD_LOOP_i_and_cse ) begin
      LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_2 <= MUX_s_1_2_2(LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_2,
          LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_1, LOAD_BATCH_LOOP_and_4_tmp);
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2 <= MUX_s_1_2_2(exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2,
          exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_1, LOAD_BATCH_LOOP_and_4_tmp);
      LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_3 <= MUX_s_1_2_2(LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_2,
          LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_3, or_dcpl_41);
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_3 <= MUX_s_1_2_2(exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2,
          exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_3, or_dcpl_41);
      exit_LOAD_BATCH_LOOP_sva_1_st_1 <= MUX1HOT_s_1_3_2((~ LOAD_BATCH_LOOP_acc_1_itm_32_1),
          exit_LOAD_BATCH_LOOP_sva_1_st, exit_LOAD_BATCH_LOOP_sva_1_st_1, {and_57_nl
          , and_58_nl , (~ LOAD_BATCH_LOOP_and_8_tmp)});
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_1 <= MUX_s_1_2_2(exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_1,
          LOAD_LOOP_LOAD_LOOP_and_cse, LOAD_BATCH_LOOP_and_8_tmp);
      LOAD_LOOP_asn_itm_1 <= MUX_s_1_2_2(LOAD_LOOP_asn_itm_1, LOAD_LOOP_asn_itm,
          LOAD_BATCH_LOOP_and_8_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_1 <= 1'b0;
    end
    else if ( LOAD_LOOP_i_and_cse & (and_dcpl_15 | and_60_rgt) ) begin
      LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm_1 <= MUX_s_1_2_2((LOAD_LOOP_acc_2_tmp[7]),
          LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm, and_60_rgt);
    end
  end
  always @(posedge clk) begin
    if ( load_wen & (~((LOAD_LOOP_acc_2_tmp[7]) | (~ LOAD_BATCH_LOOP_and_8_tmp)))
        ) begin
      LOAD_LOOP_i_7_0_lpi_1_6_0 <= LOAD_LOOP_acc_2_tmp[6:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_LOAD_BATCH_LOOP_sva_1_st <= 1'b0;
    end
    else if ( load_wen & LOAD_LOOP_asn_itm & LOAD_BATCH_LOOP_and_8_tmp ) begin
      exit_LOAD_BATCH_LOOP_sva_1_st <= ~ LOAD_BATCH_LOOP_acc_1_itm_32_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm <= 1'b0;
    end
    else if ( load_wen & (~(or_dcpl_30 | (~ (fsm_output[1])))) ) begin
      LOAD_LOOP_i_slc_LOAD_LOOP_i_7_0_7_itm <= LOAD_LOOP_acc_2_tmp[7];
    end
  end
  assign LOAD_BATCH_LOOP_b_and_nl = ((exitL_exit_LOAD_LOOP_sva & (~ LOAD_BATCH_LOOP_acc_1_itm_32_1)
      & LOAD_LOOP_asn_itm) | (LOAD_BATCH_LOOP_acc_2_tmp[4]) | (~ (LOAD_LOOP_acc_2_tmp[7]))
      | (~ LOAD_BATCH_LOOP_and_8_tmp)) & (fsm_output[1]);
  assign LOAD_BATCH_LOOP_b_mux_2_nl = MUX_v_4_2_2((LOAD_BATCH_LOOP_acc_2_tmp[3:0]),
      LOAD_BATCH_LOOP_b_4_0_sva_3_0, LOAD_BATCH_LOOP_b_and_nl);
  assign and_42_nl = and_dcpl_6 & LOAD_BATCH_LOOP_and_8_tmp & LOAD_BATCH_LOOP_stage_0;
  assign and_44_nl = (~ LOAD_BATCH_LOOP_stage_v) & LOAD_BATCH_LOOP_stage_0;
  assign or_74_nl = mux_tmp_41 | (~ LOAD_BATCH_LOOP_stage_0);
  assign LOAD_BATCH_LOOP_mux1h_nl = MUX1HOT_s_1_3_2(exitL_exit_LOAD_LOOP_sva_mx1w0,
      exitL_exit_LOAD_LOOP_sva, LOAD_LOOP_asn_itm, {and_42_nl , and_44_nl , or_74_nl});
  assign or_76_nl = LOAD_LOOP_LOAD_LOOP_and_cse | and_162_cse | (~ LOAD_BATCH_LOOP_and_8_tmp);
  assign LOAD_BATCH_LOOP_mux_26_nl = MUX_s_1_2_2(exitL_exit_LOAD_LOOP_sva_mx1w0,
      exitL_exit_LOAD_LOOP_sva, or_76_nl);
  assign LOAD_LOOP_i_nand_nl = ~((fsm_output[1]) & LOAD_BATCH_LOOP_and_8_tmp);
  assign LOAD_LOOP_i_and_4_nl = and_dcpl_56 & (fsm_output[1]);
  assign and_61_nl = (~ exitL_exit_LOAD_LOOP_sva) & LOAD_BATCH_LOOP_and_8_tmp & (fsm_output[1]);
  assign LOAD_BATCH_LOOP_mux_23_nl = MUX_s_1_2_2(LOAD_BATCH_LOOP_stage_0_1, LOAD_BATCH_LOOP_stage_0,
      LOAD_BATCH_LOOP_and_8_tmp);
  assign nor_nl = ~(LOAD_BATCH_LOOP_and_4_tmp | LOAD_BATCH_LOOP_and_8_tmp);
  assign LOAD_BATCH_LOOP_mux_25_nl = MUX_s_1_2_2(LOAD_BATCH_LOOP_stage_0_1, LOAD_BATCH_LOOP_stage_0_2,
      nor_nl);
  assign and_48_nl = or_dcpl_41 & (~ LOAD_BATCH_LOOP_and_4_tmp);
  assign LOAD_BATCH_LOOP_mux_24_nl = MUX_s_1_2_2(LOAD_BATCH_LOOP_stage_0_2, LOAD_BATCH_LOOP_stage_0_3,
      and_48_nl);
  assign and_57_nl = LOAD_LOOP_asn_itm & LOAD_BATCH_LOOP_and_8_tmp;
  assign and_58_nl = (~ LOAD_LOOP_asn_itm) & LOAD_BATCH_LOOP_and_8_tmp;

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input [0:0] vector;
  begin
    signext_7_1= {{6{vector[0]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [32:0] conv_u2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_33 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_store
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_store (
  clk, rst, conf_info, acc_done, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg,
      dma_write_chnl_val, dma_write_chnl_rdy, dma_write_chnl_msg, done, output_ready_req_req,
      output_ready_ack_ack, plm_out_cns_radr, plm_out_cns_q, plm_out_cns_req_vz,
      plm_out_cns_rls_lz
);
  input clk;
  input rst;
  input [31:0] conf_info;
  output acc_done;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;
  input done;
  input output_ready_req_req;
  output output_ready_ack_ack;
  output [6:0] plm_out_cns_radr;
  input [31:0] plm_out_cns_q;
  input plm_out_cns_req_vz;
  output plm_out_cns_rls_lz;


  // Interconnect Declarations
  wire [31:0] plm_out_cnsi_q_d;
  wire [6:0] plm_out_cnsi_radr_d;
  wire plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_softmax_sysc_store_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_7_32_128_128_32_1_gen
      plm_out_cnsi (
      .q(plm_out_cns_q),
      .radr(plm_out_cns_radr),
      .q_d(plm_out_cnsi_q_d),
      .radr_d(plm_out_cnsi_radr_d),
      .readA_r_ram_ir_internal_RMASK_B_d(plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_softmax_sysc_softmax_sysc_store_store softmax_sysc_store_store_inst (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .acc_done(acc_done),
      .dma_write_ctrl_val(dma_write_ctrl_val),
      .dma_write_ctrl_rdy(dma_write_ctrl_rdy),
      .dma_write_ctrl_msg(dma_write_ctrl_msg),
      .dma_write_chnl_val(dma_write_chnl_val),
      .dma_write_chnl_rdy(dma_write_chnl_rdy),
      .dma_write_chnl_msg(dma_write_chnl_msg),
      .done(done),
      .output_ready_req_req(output_ready_req_req),
      .output_ready_ack_ack(output_ready_ack_ack),
      .plm_out_cns_req_vz(plm_out_cns_req_vz),
      .plm_out_cns_rls_lz(plm_out_cns_rls_lz),
      .plm_out_cnsi_q_d(plm_out_cnsi_q_d),
      .plm_out_cnsi_radr_d(plm_out_cnsi_radr_d),
      .plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d(plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_compute
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_compute (
  clk, rst, conf_info, done, input_ready_req_req, input_ready_ack_ack, output_ready_req_req,
      output_ready_ack_ack, plm_in_cns_radr, plm_in_cns_q, plm_in_cns_req_vz, plm_in_cns_rls_lz,
      plm_out_cns_wadr, plm_out_cns_d, plm_out_cns_we, plm_out_cns_req_vz, plm_out_cns_rls_lz
);
  input clk;
  input rst;
  input [31:0] conf_info;
  input done;
  input input_ready_req_req;
  output input_ready_ack_ack;
  output output_ready_req_req;
  input output_ready_ack_ack;
  output [6:0] plm_in_cns_radr;
  input [31:0] plm_in_cns_q;
  input plm_in_cns_req_vz;
  output plm_in_cns_rls_lz;
  output [6:0] plm_out_cns_wadr;
  output [31:0] plm_out_cns_d;
  output plm_out_cns_we;
  input plm_out_cns_req_vz;
  output plm_out_cns_rls_lz;


  // Interconnect Declarations
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] plm_in_cnsi_q_d;
  wire [6:0] plm_in_cnsi_radr_d;
  wire plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] plm_out_cnsi_d_d;
  wire [6:0] plm_out_cnsi_wadr_d;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_clken;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_q;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_radr;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_we;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_d;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wadr;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff;
  wire plm_out_cnsi_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  BLOCK_1R1W_RBW #(.addr_width(32'sd7),
  .data_width(32'sd67),
  .depth(32'sd128),
  .latency(32'sd1)) ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_comp
      (
      .clk(clk),
      .clken(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_clken),
      .d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_d),
      .q(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_q),
      .radr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_radr),
      .wadr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wadr),
      .we(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_we)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_17_7_67_128_128_67_1_gen
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci
      (
      .clken(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_clken),
      .q(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_q),
      .radr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_radr),
      .we(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_we),
      .d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_d),
      .wadr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wadr),
      .clken_d(1'b1),
      .d_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d),
      .q_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d),
      .radr_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d),
      .wadr_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d),
      .we_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_7_32_128_128_32_1_gen
      plm_in_cnsi (
      .q(plm_in_cns_q),
      .radr(plm_in_cns_radr),
      .q_d(plm_in_cnsi_q_d),
      .radr_d(plm_in_cnsi_radr_d),
      .readA_r_ram_ir_internal_RMASK_B_d(plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_35_7_32_128_128_32_1_gen
      plm_out_cnsi (
      .we(plm_out_cns_we),
      .d(plm_out_cns_d),
      .wadr(plm_out_cns_wadr),
      .d_d(plm_out_cnsi_d_d),
      .wadr_d(plm_out_cnsi_wadr_d),
      .we_d(plm_out_cnsi_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(plm_out_cnsi_we_d_iff)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute_compute softmax_sysc_compute_compute_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .done(done),
      .input_ready_req_req(input_ready_req_req),
      .input_ready_ack_ack(input_ready_ack_ack),
      .output_ready_req_req(output_ready_req_req),
      .output_ready_ack_ack(output_ready_ack_ack),
      .plm_in_cns_req_vz(plm_in_cns_req_vz),
      .plm_in_cns_rls_lz(plm_in_cns_rls_lz),
      .plm_out_cns_req_vz(plm_out_cns_req_vz),
      .plm_out_cns_rls_lz(plm_out_cns_rls_lz),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .plm_in_cnsi_q_d(plm_in_cnsi_q_d),
      .plm_in_cnsi_radr_d(plm_in_cnsi_radr_d),
      .plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d(plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d),
      .plm_out_cnsi_d_d(plm_out_cnsi_d_d),
      .plm_out_cnsi_wadr_d(plm_out_cnsi_wadr_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff),
      .plm_out_cnsi_we_d_pff(plm_out_cnsi_we_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_load
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_load (
  clk, rst, conf_info, dma_read_ctrl_val, dma_read_ctrl_rdy, dma_read_ctrl_msg, dma_read_chnl_val,
      dma_read_chnl_rdy, dma_read_chnl_msg, done, input_ready_req_req, input_ready_ack_ack,
      plm_in_cns_wadr, plm_in_cns_d, plm_in_cns_we, plm_in_cns_req_vz, plm_in_cns_rls_lz
);
  input clk;
  input rst;
  input [31:0] conf_info;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  input done;
  output input_ready_req_req;
  input input_ready_ack_ack;
  output [6:0] plm_in_cns_wadr;
  output [31:0] plm_in_cns_d;
  output plm_in_cns_we;
  input plm_in_cns_req_vz;
  output plm_in_cns_rls_lz;


  // Interconnect Declarations
  wire [31:0] plm_in_cnsi_d_d;
  wire [6:0] plm_in_cnsi_wadr_d;
  wire plm_in_cnsi_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_softmax_sysc_load_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_33_7_32_128_128_32_1_gen
      plm_in_cnsi (
      .we(plm_in_cns_we),
      .d(plm_in_cns_d),
      .wadr(plm_in_cns_wadr),
      .d_d(plm_in_cnsi_d_d),
      .wadr_d(plm_in_cnsi_wadr_d),
      .we_d(plm_in_cnsi_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(plm_in_cnsi_we_d_iff)
    );
  esp_acc_softmax_sysc_softmax_sysc_load_load softmax_sysc_load_load_inst (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .dma_read_ctrl_val(dma_read_ctrl_val),
      .dma_read_ctrl_rdy(dma_read_ctrl_rdy),
      .dma_read_ctrl_msg(dma_read_ctrl_msg),
      .dma_read_chnl_val(dma_read_chnl_val),
      .dma_read_chnl_rdy(dma_read_chnl_rdy),
      .dma_read_chnl_msg(dma_read_chnl_msg),
      .done(done),
      .input_ready_req_req(input_ready_req_req),
      .input_ready_ack_ack(input_ready_ack_ack),
      .plm_in_cns_req_vz(plm_in_cns_req_vz),
      .plm_in_cns_rls_lz(plm_in_cns_rls_lz),
      .plm_in_cnsi_d_d(plm_in_cnsi_d_d),
      .plm_in_cnsi_wadr_d(plm_in_cnsi_wadr_d),
      .plm_in_cnsi_we_d_pff(plm_in_cnsi_we_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    softmax_sysc_acshared_fx32_dma64
// ------------------------------------------------------------------


module softmax_sysc_acshared_fx32_dma64 (
  clk, rst, conf_info, conf_done, acc_done, debug, dma_read_ctrl_val, dma_read_ctrl_rdy,
      dma_read_ctrl_msg, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg,
      dma_read_chnl_val, dma_read_chnl_rdy, dma_read_chnl_msg, dma_write_chnl_val,
      dma_write_chnl_rdy, dma_write_chnl_msg
);
  input clk;
  input rst;
  input [31:0] conf_info;
  input conf_done;
  output acc_done;
  output [31:0] debug;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;


  // Interconnect Declarations
  wire done;
  wire input_ready_req_req;
  wire input_ready_ack_ack;
  wire output_ready_req_req;
  wire output_ready_ack_ack;
  wire [6:0] plm_in_cns_wadr_nsoftmax_sysc_load_inst;
  wire [31:0] plm_in_cns_d_nsoftmax_sysc_load_inst;
  wire plm_in_cns_we_nsoftmax_sysc_load_inst;
  wire plm_in_cns_req_vz_nsoftmax_sysc_load_inst;
  wire [6:0] plm_in_cns_radr_nsoftmax_sysc_compute_inst;
  wire [31:0] plm_in_cns_q_nsoftmax_sysc_compute_inst;
  wire plm_in_cns_req_vz_nsoftmax_sysc_compute_inst;
  wire [6:0] plm_out_cns_wadr_nsoftmax_sysc_compute_inst;
  wire [31:0] plm_out_cns_d_nsoftmax_sysc_compute_inst;
  wire plm_out_cns_we_nsoftmax_sysc_compute_inst;
  wire plm_out_cns_req_vz_nsoftmax_sysc_compute_inst;
  wire plm_out_cns_we_nsoftmax_sysc_compute_inst_buz;
  wire [6:0] plm_out_cns_radr_nsoftmax_sysc_store_inst;
  wire [31:0] plm_out_cns_q_nsoftmax_sysc_store_inst;
  wire plm_out_cns_req_vz_nsoftmax_sysc_store_inst;
  wire plm_in_cns_rls_lz_nsoftmax_sysc_load_inst_bud;
  wire plm_in_cns_rls_lz_nsoftmax_sysc_compute_inst_bud;
  wire plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud;
  wire plm_out_cns_rls_lz_nsoftmax_sysc_compute_inst_bud;
  wire plm_out_cns_rls_lz_nsoftmax_sysc_store_inst_bud;
  wire plm_in_cns_R0;
  wire plm_in_cns_S1;
  wire plm_in_cns_R1;
  wire [31:0] plm_in_cns_d_shi0;
  wire [31:0] plm_in_cns_d_shi1;
  wire [31:0] plm_in_cns_q_sho0;
  wire [31:0] plm_in_cns_q_sho1;
  wire [6:0] plm_in_cns_radr_shi0;
  wire [6:0] plm_in_cns_radr_shi1;
  wire [6:0] plm_in_cns_wadr_shi0;
  wire [6:0] plm_in_cns_wadr_shi1;
  wire plm_in_cns_we_shi0;
  wire plm_in_cns_we_shi1;
  wire plm_out_cns_R0;
  wire plm_out_cns_S1;
  wire plm_out_cns_R1;
  wire [31:0] plm_out_cns_d_shi0;
  wire [31:0] plm_out_cns_d_shi1;
  wire [31:0] plm_out_cns_q_sho0;
  wire [31:0] plm_out_cns_q_sho1;
  wire [6:0] plm_out_cns_radr_shi0;
  wire [6:0] plm_out_cns_radr_shi1;
  wire [6:0] plm_out_cns_wadr_shi0;
  wire [6:0] plm_out_cns_wadr_shi1;
  wire plm_out_cns_we_shi0;
  wire plm_out_cns_we_shi1;
  wire plm_in_cns_S0_iff;
  wire plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_iff;
  wire plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud_iff;
  wire plm_out_cns_S0_iff;
  wire plm_in_cns_S0_dmo;
  wire plm_out_cns_S0_dmo;


  // Interconnect Declarations for Component Instantiations 
  BLOCK_1R1W_RBW #(.addr_width(32'sd7),
  .data_width(32'sd32),
  .depth(32'sd128),
  .latency(32'sd1)) plm_in_cns_comp (
      .clk(clk),
      .clken(1'b1),
      .d(plm_in_cns_d_shi0),
      .q(plm_in_cns_q_sho0),
      .radr(plm_in_cns_radr_shi0),
      .wadr(plm_in_cns_wadr_shi0),
      .we(plm_in_cns_we_shi0)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd7),
  .data_width(32'sd32),
  .depth(32'sd128),
  .latency(32'sd1)) plm_in_cns_comp_1 (
      .clk(clk),
      .clken(1'b1),
      .d(plm_in_cns_d_shi1),
      .q(plm_in_cns_q_sho1),
      .radr(plm_in_cns_radr_shi1),
      .wadr(plm_in_cns_wadr_shi1),
      .we(plm_in_cns_we_shi1)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd7),
  .data_width(32'sd32),
  .depth(32'sd128),
  .latency(32'sd1)) plm_out_cns_comp (
      .clk(clk),
      .clken(1'b1),
      .d(plm_out_cns_d_shi0),
      .q(plm_out_cns_q_sho0),
      .radr(plm_out_cns_radr_shi0),
      .wadr(plm_out_cns_wadr_shi0),
      .we(plm_out_cns_we_shi0)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd7),
  .data_width(32'sd32),
  .depth(32'sd128),
  .latency(32'sd1)) plm_out_cns_comp_1 (
      .clk(clk),
      .clken(1'b1),
      .d(plm_out_cns_d_shi1),
      .q(plm_out_cns_q_sho1),
      .radr(plm_out_cns_radr_shi1),
      .wadr(plm_out_cns_wadr_shi1),
      .we(plm_out_cns_we_shi1)
    );
  esp_acc_softmax_sysc_softmax_sysc_load softmax_sysc_load_inst (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .dma_read_ctrl_val(dma_read_ctrl_val),
      .dma_read_ctrl_rdy(dma_read_ctrl_rdy),
      .dma_read_ctrl_msg(dma_read_ctrl_msg),
      .dma_read_chnl_val(dma_read_chnl_val),
      .dma_read_chnl_rdy(dma_read_chnl_rdy),
      .dma_read_chnl_msg(dma_read_chnl_msg),
      .done(done),
      .input_ready_req_req(input_ready_req_req),
      .input_ready_ack_ack(input_ready_ack_ack),
      .plm_in_cns_wadr(plm_in_cns_wadr_nsoftmax_sysc_load_inst),
      .plm_in_cns_d(plm_in_cns_d_nsoftmax_sysc_load_inst),
      .plm_in_cns_we(plm_in_cns_we_nsoftmax_sysc_load_inst),
      .plm_in_cns_req_vz(plm_in_cns_req_vz_nsoftmax_sysc_load_inst),
      .plm_in_cns_rls_lz(plm_in_cns_rls_lz_nsoftmax_sysc_load_inst_bud)
    );
  esp_acc_softmax_sysc_softmax_sysc_compute softmax_sysc_compute_inst (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .done(done),
      .input_ready_req_req(input_ready_req_req),
      .input_ready_ack_ack(input_ready_ack_ack),
      .output_ready_req_req(output_ready_req_req),
      .output_ready_ack_ack(output_ready_ack_ack),
      .plm_in_cns_radr(plm_in_cns_radr_nsoftmax_sysc_compute_inst),
      .plm_in_cns_q(plm_in_cns_q_nsoftmax_sysc_compute_inst),
      .plm_in_cns_req_vz(plm_in_cns_req_vz_nsoftmax_sysc_compute_inst),
      .plm_in_cns_rls_lz(plm_in_cns_rls_lz_nsoftmax_sysc_compute_inst_bud),
      .plm_out_cns_wadr(plm_out_cns_wadr_nsoftmax_sysc_compute_inst),
      .plm_out_cns_d(plm_out_cns_d_nsoftmax_sysc_compute_inst),
      .plm_out_cns_we(plm_out_cns_we_nsoftmax_sysc_compute_inst),
      .plm_out_cns_req_vz(plm_out_cns_req_vz_nsoftmax_sysc_compute_inst),
      .plm_out_cns_rls_lz(plm_out_cns_rls_lz_nsoftmax_sysc_compute_inst_bud)
    );
  esp_acc_softmax_sysc_softmax_sysc_store softmax_sysc_store_inst (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .acc_done(acc_done),
      .dma_write_ctrl_val(dma_write_ctrl_val),
      .dma_write_ctrl_rdy(dma_write_ctrl_rdy),
      .dma_write_ctrl_msg(dma_write_ctrl_msg),
      .dma_write_chnl_val(dma_write_chnl_val),
      .dma_write_chnl_rdy(dma_write_chnl_rdy),
      .dma_write_chnl_msg(dma_write_chnl_msg),
      .done(done),
      .output_ready_req_req(output_ready_req_req),
      .output_ready_ack_ack(output_ready_ack_ack),
      .plm_out_cns_radr(plm_out_cns_radr_nsoftmax_sysc_store_inst),
      .plm_out_cns_q(plm_out_cns_q_nsoftmax_sysc_store_inst),
      .plm_out_cns_req_vz(plm_out_cns_req_vz_nsoftmax_sysc_store_inst),
      .plm_out_cns_rls_lz(plm_out_cns_rls_lz_nsoftmax_sysc_store_inst_bud)
    );
  esp_acc_softmax_sysc_unreg_hier unreg (
      .in_0(plm_in_cns_S0_iff),
      .out_0(plm_in_cns_R0)
    );
  esp_acc_softmax_sysc_unreg_hier unreg_1 (
      .in_0(plm_in_cns_S1),
      .out_0(plm_in_cns_R1)
    );
  esp_acc_softmax_sysc_unreg_hier unreg_2 (
      .in_0(plm_out_cns_S0_iff),
      .out_0(plm_out_cns_R0)
    );
  esp_acc_softmax_sysc_unreg_hier unreg_3 (
      .in_0(plm_out_cns_S1),
      .out_0(plm_out_cns_R1)
    );
  esp_acc_softmax_sysc_softmax_sysc_plm_in_cns_bctl softmax_sysc_plm_in_cns_bctl_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_wadr_nsoftmax_sysc_load_inst(plm_in_cns_wadr_nsoftmax_sysc_load_inst),
      .plm_in_cns_d_nsoftmax_sysc_load_inst(plm_in_cns_d_nsoftmax_sysc_load_inst),
      .plm_in_cns_we_nsoftmax_sysc_load_inst(plm_in_cns_we_nsoftmax_sysc_load_inst),
      .plm_in_cns_req_vz_nsoftmax_sysc_load_inst(plm_in_cns_req_vz_nsoftmax_sysc_load_inst),
      .plm_in_cns_radr_nsoftmax_sysc_compute_inst(plm_in_cns_radr_nsoftmax_sysc_compute_inst),
      .plm_in_cns_q_nsoftmax_sysc_compute_inst(plm_in_cns_q_nsoftmax_sysc_compute_inst),
      .plm_in_cns_req_vz_nsoftmax_sysc_compute_inst(plm_in_cns_req_vz_nsoftmax_sysc_compute_inst),
      .plm_out_cns_we_nsoftmax_sysc_compute_inst_buz(plm_out_cns_we_nsoftmax_sysc_compute_inst_buz),
      .plm_in_cns_rls_lz_nsoftmax_sysc_load_inst_bud(plm_in_cns_rls_lz_nsoftmax_sysc_load_inst_bud),
      .plm_in_cns_rls_lz_nsoftmax_sysc_compute_inst_bud(plm_in_cns_rls_lz_nsoftmax_sysc_compute_inst_bud),
      .plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud(plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud),
      .plm_out_cns_rls_lz_nsoftmax_sysc_compute_inst_bud(1'b0),
      .plm_in_cns_S0(plm_in_cns_S0_dmo),
      .plm_in_cns_R0(plm_in_cns_R0),
      .plm_in_cns_S1(plm_in_cns_S1),
      .plm_in_cns_R1(plm_in_cns_R1),
      .plm_in_cns_d_shi0(plm_in_cns_d_shi0),
      .plm_in_cns_d_shi1(plm_in_cns_d_shi1),
      .plm_in_cns_q_sho0(plm_in_cns_q_sho0),
      .plm_in_cns_q_sho1(plm_in_cns_q_sho1),
      .plm_in_cns_radr_shi0(plm_in_cns_radr_shi0),
      .plm_in_cns_radr_shi1(plm_in_cns_radr_shi1),
      .plm_in_cns_wadr_shi0(plm_in_cns_wadr_shi0),
      .plm_in_cns_wadr_shi1(plm_in_cns_wadr_shi1),
      .plm_in_cns_we_shi0(plm_in_cns_we_shi0),
      .plm_in_cns_we_shi1(plm_in_cns_we_shi1),
      .plm_in_cns_S0_pff(plm_in_cns_S0_iff),
      .plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_pff(plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_iff),
      .plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud_pff(plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud_iff)
    );
  esp_acc_softmax_sysc_softmax_sysczjlBRut_cns_bctl softmax_sysczjlBRut_cns_bctl_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_wadr_nsoftmax_sysc_compute_inst(plm_out_cns_wadr_nsoftmax_sysc_compute_inst),
      .plm_out_cns_d_nsoftmax_sysc_compute_inst(plm_out_cns_d_nsoftmax_sysc_compute_inst),
      .plm_out_cns_we_nsoftmax_sysc_compute_inst(plm_out_cns_we_nsoftmax_sysc_compute_inst),
      .plm_out_cns_req_vz_nsoftmax_sysc_compute_inst(plm_out_cns_req_vz_nsoftmax_sysc_compute_inst),
      .plm_out_cns_we_nsoftmax_sysc_compute_inst_buz(1'b0),
      .plm_out_cns_radr_nsoftmax_sysc_store_inst(plm_out_cns_radr_nsoftmax_sysc_store_inst),
      .plm_out_cns_q_nsoftmax_sysc_store_inst(plm_out_cns_q_nsoftmax_sysc_store_inst),
      .plm_out_cns_req_vz_nsoftmax_sysc_store_inst(plm_out_cns_req_vz_nsoftmax_sysc_store_inst),
      .plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud(plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud),
      .plm_out_cns_rls_lz_nsoftmax_sysc_compute_inst_bud(plm_out_cns_rls_lz_nsoftmax_sysc_compute_inst_bud),
      .plm_out_cns_rls_lz_nsoftmax_sysc_store_inst_bud(plm_out_cns_rls_lz_nsoftmax_sysc_store_inst_bud),
      .plm_out_cns_S0(plm_out_cns_S0_dmo),
      .plm_out_cns_R0(plm_out_cns_R0),
      .plm_out_cns_S1(plm_out_cns_S1),
      .plm_out_cns_R1(plm_out_cns_R1),
      .plm_out_cns_d_shi0(plm_out_cns_d_shi0),
      .plm_out_cns_d_shi1(plm_out_cns_d_shi1),
      .plm_out_cns_q_sho0(plm_out_cns_q_sho0),
      .plm_out_cns_q_sho1(plm_out_cns_q_sho1),
      .plm_out_cns_radr_shi0(plm_out_cns_radr_shi0),
      .plm_out_cns_radr_shi1(plm_out_cns_radr_shi1),
      .plm_out_cns_wadr_shi0(plm_out_cns_wadr_shi0),
      .plm_out_cns_wadr_shi1(plm_out_cns_wadr_shi1),
      .plm_out_cns_we_shi0(plm_out_cns_we_shi0),
      .plm_out_cns_we_shi1(plm_out_cns_we_shi1),
      .plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_pff(plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_iff),
      .plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud_pff(plm_out_cns_we_nsoftmax_sysc_compute_inst_buz_bud_iff),
      .plm_out_cns_S0_pff(plm_out_cns_S0_iff)
    );
  esp_acc_softmax_sysc_softmax_sysc_config softmax_sysc_config_inst (
      .clk(clk),
      .rst(rst),
      .conf_done(conf_done),
      .done(done)
    );
  assign debug = 32'b00000000000000000000000000000000;
endmodule



