
//------> ./softmax_Connections_OutBlockingless_dma_info_tcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_Connections_OutBlockingless_dma_info_tcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_Connections_OutBlockingless_dma_info_tcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue May 19 12:17:59 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core
    (
  this_val, this_rdy, this_msg, m_index_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [66:0] this_msg;
  input [31:0] m_index_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire [31:0] m_index_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [24:0] m_index_slc_m_index_31_7_psp_lpi_1_dfm;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  reg reg_128_3_reg_7;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd32)) m_index_rsci (
      .dat(m_index_rsc_dat),
      .idat(m_index_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd45),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 #(.rscid(32'sd50)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign this_msg = {27'b000000000000000000000000000 , reg_128_3_reg_7 , 7'b0000000
      , m_index_slc_m_index_31_7_psp_lpi_1_dfm , 7'b0000000};
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      reg_128_3_reg_7 <= 1'b0;
    end
    else if ( (~((~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1) | this_rdy)) | ccs_ccore_start_rsci_idat
        ) begin
      reg_128_3_reg_7 <= 1'b1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_val <= 1'b0;
    end
    else if ( or_4_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      m_index_slc_m_index_31_7_psp_lpi_1_dfm <= 25'b0000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      m_index_slc_m_index_31_7_psp_lpi_1_dfm <= m_index_rsci_idat[31:7];
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module esp_acc_softmax_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_index_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  input this_rdy;
  output [66:0] this_msg;
  input [31:0] m_index_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_esp_acc_softmax_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core_inst (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_index_rsc_dat(m_index_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_Connections_InBlockingless_sc_dt_sc_bvless_64greater_comma_Connections_SYN_PORTgreater_Pop_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./softmax_Connections_InBlockingless_sc_dt_sc_bvless_64greater_comma_Connections_SYN_PORTgreater_Pop_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_Connections_InBlockingless_sc_dt_sc_bvless_64greater_comma_Connections_SYN_PORTgreater_Pop_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_Connections_InBlockingless_sc_dt_sc_bvless_64greater_comma_Connections_SYN_PORTgreater_Pop.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue May 19 11:53:49 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_Connections_InBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Pop_core
// ------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_Connections_InBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Pop_core
    (
  this_val, this_rdy, this_msg, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [63:0] this_msg;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_2_cse;
  wire this_rdy_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [63:0] nl_return_rsci_d;
  assign nl_return_rsci_d = this_msg;
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_val;
  esp_acc_softmax_esp_acc_softmax_mgc_out_dreg_v2 #(.rscid(32'sd4),
  .width(32'sd64)) return_rsci (
      .d(nl_return_rsci_d[63:0]),
      .z(return_rsc_z)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd44),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 #(.rscid(32'sd49)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign or_2_cse = ccs_ccore_start_rsci_idat | (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_val));
  assign this_rdy_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_val
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_rdy <= 1'b0;
    end
    else if ( or_2_cse | this_rdy_mx0c1 ) begin
      this_rdy <= ~ this_rdy_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_2_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Pop
// ------------------------------------------------------------------


module esp_acc_softmax_Connections_InBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Pop (
  this_val, this_rdy, this_msg, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  input this_val;
  output this_rdy;
  input [63:0] this_msg;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_esp_acc_softmax_Connections_InBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Pop_core
      Connections_InBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Pop_core_inst (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_handshake_t_req_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_handshake_t_req_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_handshake_t_req.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue May 19 11:53:48 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_handshake_t_req_core
// ------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_handshake_t_req_core (
  this_req_req, this_ack_ack, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld, ccs_MIO_clk,
      ccs_MIO_srst
);
  output this_req_req;
  reg this_req_req;
  input this_ack_ack;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg do_asn_mdf_sva_st_1;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_st_2;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = do_asn_mdf_sva_st_1 & io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_st_2;
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd43),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 #(.rscid(32'sd48)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_req_req <= 1'b0;
      do_asn_mdf_sva_st_1 <= 1'b0;
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_st_2 <= 1'b0;
    end
    else begin
      this_req_req <= io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_ack_ack;
      do_asn_mdf_sva_st_1 <= this_ack_ack;
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= ccs_ccore_start_rsci_idat |
          (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_ack_ack));
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_st_2 <= io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    handshake_t_req
// ------------------------------------------------------------------


module esp_acc_softmax_handshake_t_req (
  this_req_req, this_ack_ack, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld, ccs_MIO_clk,
      ccs_MIO_srst
);
  output this_req_req;
  input this_ack_ack;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_esp_acc_softmax_handshake_t_req_core handshake_t_req_core_inst (
      .this_req_req(this_req_req),
      .this_ack_ack(this_ack_ack),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./softmax_mgc_in_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_mgc_in_sync_v2 (vd, vz);
    parameter valid = 1;

    output vd;
    input  vz;

    wire   vd;

    assign vd = vz;

endmodule



//------> ./softmax_handshake_t_ack_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_handshake_t_ack_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_handshake_t_ack.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue May 19 11:53:47 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_handshake_t_ack_core
// ------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_handshake_t_ack_core (
  this_req_req, this_ack_ack, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld, ccs_MIO_clk,
      ccs_MIO_srst
);
  input this_req_req;
  output this_ack_ack;
  reg this_ack_ack;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire asn_ccs_ccore_done_synci_ivld_and_cse;
  wire this_ack_ack_mx0c1;


  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd42),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 #(.rscid(32'sd47)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(asn_ccs_ccore_done_synci_ivld_and_cse)
    );
  assign asn_ccs_ccore_done_synci_ivld_and_cse = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_req_req;
  assign this_ack_ack_mx0c1 = asn_ccs_ccore_done_synci_ivld_and_cse & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_ack_ack <= 1'b0;
    end
    else if ( (((~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1) | this_req_req) &
        ccs_ccore_start_rsci_idat) | this_ack_ack_mx0c1 ) begin
      this_ack_ack <= ~ this_ack_ack_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( ~(io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_req_req)) )
        begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    handshake_t_ack
// ------------------------------------------------------------------


module esp_acc_softmax_handshake_t_ack (
  this_req_req, this_ack_ack, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld, ccs_MIO_clk,
      ccs_MIO_srst
);
  input this_req_req;
  output this_ack_ack;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_esp_acc_softmax_handshake_t_ack_core handshake_t_ack_core_inst (
      .this_req_req(this_req_req),
      .this_ack_ack(this_ack_ack),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_mgc_shift_br_beh_v5.v 
module esp_acc_softmax_mgc_shift_br_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_s(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_s(a,s,1'b0);
     end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshr_u

   //Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction

endmodule

//------> ./softmax_mgc_shift_bl_beh_v5.v 
module esp_acc_softmax_mgc_shift_bl_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate if ( signd_a )
   begin: SGNED
     assign z = fshl_s(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
     assign z = fshl_s(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

endmodule

//------> ./softmax_mgc_shift_l_beh_v5.v 
module esp_acc_softmax_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./softmax_leading_sign_74_0.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Wed Apr 29 22:59:54 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_74_0
// ------------------------------------------------------------------


module esp_acc_softmax_leading_sign_74_0 (
  mantissa, rtn
);
  input [73:0] mantissa;
  output [6:0] rtn;


  // Interconnect Declarations
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_24;
  wire c_h_1_27;
  wire c_h_1_28;
  wire c_h_1_29;
  wire c_h_1_30;
  wire c_h_1_33;
  wire c_h_1_34;
  wire c_h_1_35;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc;

  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_1_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_292_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_2_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_or_2_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_nor_nl;

  // Interconnect Declarations for Component Instantiations
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2
      = ~((mantissa[71:70]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1
      = ~((mantissa[73:72]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1
      = ~((mantissa[69:68]!=2'b00));
  assign c_h_1_2 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3
      = (mantissa[67:66]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2
      = ~((mantissa[63:62]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1
      = ~((mantissa[65:64]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1
      = ~((mantissa[61:60]!=2'b00));
  assign c_h_1_5 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4
      = (mantissa[59:58]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1
      & c_h_1_5;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2
      = ~((mantissa[55:54]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1
      = ~((mantissa[57:56]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1
      = ~((mantissa[53:52]!=2'b00));
  assign c_h_1_9 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3
      = (mantissa[51:50]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2
      = ~((mantissa[47:46]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1
      = ~((mantissa[49:48]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1
      = ~((mantissa[45:44]!=2'b00));
  assign c_h_1_12 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5
      = (mantissa[43:42]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1
      & c_h_1_12 & c_h_1_13;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2
      = ~((mantissa[39:38]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1
      = ~((mantissa[41:40]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1
      = ~((mantissa[37:36]!=2'b00));
  assign c_h_1_17 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3
      = (mantissa[35:34]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2
      = ~((mantissa[31:30]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1
      = ~((mantissa[33:32]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1
      = ~((mantissa[29:28]!=2'b00));
  assign c_h_1_20 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4
      = (mantissa[27:26]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1
      & c_h_1_20;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2
      = ~((mantissa[23:22]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1
      = ~((mantissa[25:24]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1
      = ~((mantissa[21:20]!=2'b00));
  assign c_h_1_24 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3
      = (mantissa[19:18]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2
      = ~((mantissa[15:14]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1
      = ~((mantissa[17:16]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1
      = ~((mantissa[13:12]!=2'b00));
  assign c_h_1_27 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2;
  assign c_h_1_28 = c_h_1_24 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3;
  assign c_h_1_29 = c_h_1_21 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_30 = c_h_1_14 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6
      = (mantissa[11:10]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1
      & c_h_1_27 & c_h_1_28 & c_h_1_29;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2
      = ~((mantissa[7:6]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1
      = ~((mantissa[9:8]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1
      = ~((mantissa[5:4]!=2'b00));
  assign c_h_1_33 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3
      = (mantissa[3:2]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1;
  assign c_h_1_34 = c_h_1_33 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3;
  assign c_h_1_35 = c_h_1_30 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc
      = (mantissa[1:0]==2'b00) & c_h_1_34 & c_h_1_35;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_nl
      = c_h_1_30 & (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6);
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_1_nl
      = c_h_1_14 & (c_h_1_29 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5))
      & (~ c_h_1_35);
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_292_nl
      = c_h_1_6 & (c_h_1_13 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4))
      & (~((~(c_h_1_21 & (c_h_1_28 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4))))
      & c_h_1_30)) & (c_h_1_34 | (~ c_h_1_35));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_2_nl
      = c_h_1_2 & (c_h_1_5 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3))
      & (~((~(c_h_1_9 & (c_h_1_12 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~((~(c_h_1_17 & (c_h_1_20 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3))
      & (~((~(c_h_1_24 & (c_h_1_27 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3))))
      & c_h_1_29)))) & c_h_1_30)) & (~((~(c_h_1_33 & (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3)))
      & c_h_1_35));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_or_2_nl
      = (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2))))
      & c_h_1_21)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2))))
      & c_h_1_28)))) & c_h_1_29)))) & c_h_1_30)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2))
      & (~ c_h_1_34))) & c_h_1_35))) | ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_nor_nl
      = ~((mantissa[73]) | (~((mantissa[72:71]!=2'b01))) | (((mantissa[69]) | (~((mantissa[68:67]!=2'b01))))
      & c_h_1_2) | ((~((~((mantissa[65]) | (~((mantissa[64:63]!=2'b01))))) & (~(((mantissa[61])
      | (~((mantissa[60:59]!=2'b01)))) & c_h_1_5)))) & c_h_1_6) | ((~((~((mantissa[57])
      | (~((mantissa[56:55]!=2'b01))))) & (~(((mantissa[53]) | (~((mantissa[52:51]!=2'b01))))
      & c_h_1_9)) & (~((~((~((mantissa[49]) | (~((mantissa[48:47]!=2'b01))))) & (~(((mantissa[45])
      | (~((mantissa[44:43]!=2'b01)))) & c_h_1_12)))) & c_h_1_13)))) & c_h_1_14)
      | ((~((~((mantissa[41]) | (~((mantissa[40:39]!=2'b01))))) & (~(((mantissa[37])
      | (~((mantissa[36:35]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[33]) | (~((mantissa[32:31]!=2'b01)))))
      & (~(((mantissa[29]) | (~((mantissa[28:27]!=2'b01)))) & c_h_1_20)))) & c_h_1_21))
      & (~((~((~((mantissa[25]) | (~((mantissa[24:23]!=2'b01))))) & (~(((mantissa[21])
      | (~((mantissa[20:19]!=2'b01)))) & c_h_1_24)) & (~((~((~((mantissa[17]) | (~((mantissa[16:15]!=2'b01)))))
      & (~(((mantissa[13]) | (~((mantissa[12:11]!=2'b01)))) & c_h_1_27)))) & c_h_1_28))))
      & c_h_1_29)))) & c_h_1_30) | ((~((~((mantissa[9]) | (~((mantissa[8:7]!=2'b01)))))
      & (~(((mantissa[5]) | (~((mantissa[4:3]!=2'b01)))) & c_h_1_33)) & (~((mantissa[1])
      & c_h_1_34)))) & c_h_1_35) | ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc);
  assign rtn = {c_h_1_35 , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_1_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_292_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_2_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_or_2_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_nor_nl};
endmodule




//------> ./softmax_mgc_mul_pipe_beh.v 
//
// File:      $Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v
//
// BASELINE:  Catapult-C version 2006b.63
// MODIFIED:  2007-04-03, tnagler
//
// Note: this file uses Verilog2001 features;
//       please enable Verilog2001 in the flow!

module esp_acc_softmax_mgc_mul_pipe (a, b, clk, en, a_rst, s_rst, z);

    // Parameters:
    parameter integer width_a = 32'd4;  // input a bit width
    parameter         signd_a =  1'b1;  // input a type (1=signed, 0=unsigned)
    parameter integer width_b = 32'd4;  // input b bit width
    parameter         signd_b =  1'b1;  // input b type (1=signed, 0=unsigned)
    parameter integer width_z = 32'd8;  // result bit width (= width_a + width_b)
    parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
    parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
    parameter    a_rst_active =  1'b1;  // unused
    parameter    s_rst_active =  1'b1;  // unused
    parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
    parameter integer n_inreg = 32'd0;  // number of input registers

    localparam integer width_ab = width_a + width_b;  // multiplier result width
    localparam integer n_inreg_min = (n_inreg > 1) ? (n_inreg-1) : 0; // for Synopsys DC

    // I/O ports:
    input  [width_a-1:0] a;      // input A
    input  [width_b-1:0] b;      // input B
    input                clk;    // clock
    input                en;     // enable
    input                a_rst;  // async reset (unused)
    input                s_rst;  // sync reset (unused)
    output [width_z-1:0] z;      // output


    // Input registers:

    wire [width_a-1:0] a_f;
    wire [width_b-1:0] b_f;

    integer i;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(negedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i];
                    b_reg[i+1] <= b_reg[i];
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    else
    begin: POS_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(posedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i];
                    b_reg[i+1] <= b_reg[i];
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    endgenerate


    // Output:
    wire [width_z-1:0]  xz;

    function signed [width_z-1:0] conv_signed;
      input signed [width_ab-1:0] res;
      conv_signed = res[width_z-1:0];
    endfunction

    generate
      wire signed [width_ab-1:0] res;
      if ( (signd_a == 1'b1) && (signd_b == 1'b1) )
      begin: SIGNED_AB
              assign res = $signed(a_f) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b1) && (signd_b == 1'b0) )
      begin: SIGNED_A
              assign res = $signed(a_f) * $signed({1'b0, b_f});
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b0) && (signd_b == 1'b1) )
      begin: SIGNED_B
              assign res = $signed({1'b0,a_f}) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else
      begin: UNSIGNED_AB
              assign res = a_f * b_f;
	      assign xz = res[width_z-1:0];
      end
    endgenerate


    // Output registers:

    reg  [width_z-1:0] reg_array[stages-2:0];
    wire [width_z-1:0] z;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE2
        always @(negedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz;
                else
                    reg_array[i] <= reg_array[i-1];
    end
    else
    begin: POS_EDGE2
        always @(posedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz;
                else
                    reg_array[i] <= reg_array[i-1];
    end
    endgenerate

    assign z = reg_array[stages-2];
endmodule

//------> /opt/cad/catapult/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 
  
)( clk,clken,d,q,radr,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" *)
  reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block"
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./softmax_Connections_OutBlockingless_sc_dt_sc_bvless_64greater_comma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_Connections_OutBlockingless_sc_dt_sc_bvless_64greater_comma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_Connections_OutBlockingless_sc_dt_sc_bvless_64greater_comma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue May 19 11:53:44 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_Connections_OutBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_Connections_OutBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Push_core
    (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [63:0] this_msg;
  input [63:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire [63:0] m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [31:0] m_slc_m_31_0_psp_lpi_1_dfm;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  reg reg_C_32_11011110101011011011111011101111_1_reg_30;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd64)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd41),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 #(.rscid(32'sd46)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign this_msg = signext_64_63({reg_C_32_11011110101011011011111011101111_1_reg_30
      , 1'b0 , ({{3{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , reg_C_32_11011110101011011011111011101111_1_reg_30 , 1'b0 , reg_C_32_11011110101011011011111011101111_1_reg_30
      , 1'b0 , ({{1{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{1{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{4{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{2{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{3{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , m_slc_m_31_0_psp_lpi_1_dfm});
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_val <= 1'b0;
    end
    else if ( or_4_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      reg_C_32_11011110101011011011111011101111_1_reg_30 <= 1'b0;
    end
    else if ( (~((~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1) | this_rdy)) | ccs_ccore_start_rsci_idat
        ) begin
      reg_C_32_11011110101011011011111011101111_1_reg_30 <= 1'b1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      m_slc_m_31_0_psp_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      m_slc_m_31_0_psp_lpi_1_dfm <= m_rsci_idat[31:0];
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end

  function automatic [63:0] signext_64_63;
    input [62:0] vector;
  begin
    signext_64_63= {{1{vector[62]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module esp_acc_softmax_Connections_OutBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  input this_rdy;
  output [63:0] this_msg;
  input [63:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_esp_acc_softmax_Connections_OutBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Push_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_rsc_dat(m_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue May 19 12:18:18 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_plm_out_cns_bctl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_plm_out_cns_bctl (
  clk, rst, plm_out_cns_wadr_nsoftmax_compute_kernel_inst, plm_out_cns_d_nsoftmax_compute_kernel_inst,
      plm_out_cns_we_nsoftmax_compute_kernel_inst, plm_out_cns_req_vz_nsoftmax_compute_kernel_inst,
      plm_out_cns_we_nsoftmax_compute_kernel_inst_buz, plm_out_cns_radr_nsoftmax_store_output_inst,
      plm_out_cns_q_nsoftmax_store_output_inst, plm_out_cns_req_vz_nsoftmax_store_output_inst,
      plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud, plm_out_cns_rls_lz_nsoftmax_compute_kernel_inst_bud,
      plm_out_cns_rls_lz_nsoftmax_store_output_inst_bud, plm_out_cns_S0, plm_out_cns_R0,
      plm_out_cns_S1, plm_out_cns_R1, plm_out_cns_d_shi0, plm_out_cns_d_shi1, plm_out_cns_q_sho0,
      plm_out_cns_q_sho1, plm_out_cns_radr_shi0, plm_out_cns_radr_shi1, plm_out_cns_wadr_shi0,
      plm_out_cns_wadr_shi1, plm_out_cns_we_shi0, plm_out_cns_we_shi1, plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_pff,
      plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud_pff, plm_out_cns_S0_pff
);
  input clk;
  input rst;
  input [6:0] plm_out_cns_wadr_nsoftmax_compute_kernel_inst;
  input [31:0] plm_out_cns_d_nsoftmax_compute_kernel_inst;
  input plm_out_cns_we_nsoftmax_compute_kernel_inst;
  output plm_out_cns_req_vz_nsoftmax_compute_kernel_inst;
  input plm_out_cns_we_nsoftmax_compute_kernel_inst_buz;
  input [6:0] plm_out_cns_radr_nsoftmax_store_output_inst;
  output [31:0] plm_out_cns_q_nsoftmax_store_output_inst;
  output plm_out_cns_req_vz_nsoftmax_store_output_inst;
  output plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud;
  input plm_out_cns_rls_lz_nsoftmax_compute_kernel_inst_bud;
  input plm_out_cns_rls_lz_nsoftmax_store_output_inst_bud;
  output plm_out_cns_S0;
  input plm_out_cns_R0;
  output plm_out_cns_S1;
  input plm_out_cns_R1;
  output [31:0] plm_out_cns_d_shi0;
  output [31:0] plm_out_cns_d_shi1;
  input [31:0] plm_out_cns_q_sho0;
  input [31:0] plm_out_cns_q_sho1;
  output [6:0] plm_out_cns_radr_shi0;
  output [6:0] plm_out_cns_radr_shi1;
  output [6:0] plm_out_cns_wadr_shi0;
  output [6:0] plm_out_cns_wadr_shi1;
  output plm_out_cns_we_shi0;
  output plm_out_cns_we_shi1;
  input plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_pff;
  output plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud_pff;
  output plm_out_cns_S0_pff;


  // Interconnect Declarations
  reg plm_out_cns_we_nsoftmax_compute_kernel_inst_buy;
  wire plm_out_cns_PC0;
  reg plm_out_cns_ppidx;
  reg [1:0] plm_out_cns_ppown;
  wire plm_out_cns_PC1;
  reg plm_out_cns_ppidx_1;
  reg [1:0] plm_out_cns_ppown_1;
  wire [1:0] plm_out_acc_rmff;
  wire [3:0] nl_plm_out_acc_rmff;
  wire plm_out_xor_rmff;
  wire [1:0] plm_out_acc_1_rmff;
  wire [3:0] nl_plm_out_acc_1_rmff;


  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_req_vz_nsoftmax_compute_kernel_inst = plm_out_cns_R0;
  assign plm_out_cns_req_vz_nsoftmax_store_output_inst = plm_out_cns_R1;
  assign plm_out_xor_rmff = plm_out_cns_ppidx ^ plm_out_cns_PC0;
  assign nl_plm_out_acc_rmff = plm_out_cns_ppown + conv_u2u_1_2(plm_out_cns_PC0)
      + conv_s2u_1_2(plm_out_cns_PC1);
  assign plm_out_acc_rmff = nl_plm_out_acc_rmff[1:0];
  assign plm_out_cns_PC0 = plm_out_cns_S0 & plm_out_cns_rls_lz_nsoftmax_compute_kernel_inst_bud;
  assign nl_plm_out_acc_1_rmff = plm_out_cns_ppown_1 + conv_u2u_1_2(plm_out_cns_PC1)
      + conv_s2u_1_2(plm_out_cns_PC0);
  assign plm_out_acc_1_rmff = nl_plm_out_acc_1_rmff[1:0];
  assign plm_out_cns_PC1 = ((plm_out_cns_ppown_1!=2'b00)) & plm_out_cns_rls_lz_nsoftmax_store_output_inst_bud;
  assign plm_out_cns_q_nsoftmax_store_output_inst = MUX_v_32_2_2(plm_out_cns_q_sho0,
      plm_out_cns_q_sho1, plm_out_cns_ppidx_1);
  assign plm_out_cns_d_shi0 = plm_out_cns_d_nsoftmax_compute_kernel_inst;
  assign plm_out_cns_radr_shi0 = plm_out_cns_radr_nsoftmax_store_output_inst;
  assign plm_out_cns_wadr_shi0 = plm_out_cns_wadr_nsoftmax_compute_kernel_inst;
  assign plm_out_cns_we_shi0 = plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_pff
      & plm_out_cns_S0_pff & (~ plm_out_xor_rmff);
  assign plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud = plm_out_cns_we_nsoftmax_compute_kernel_inst_buy;
  assign plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud_pff = plm_out_cns_we_nsoftmax_compute_kernel_inst;
  assign plm_out_cns_S0 = ~((plm_out_cns_ppown==2'b10));
  assign plm_out_cns_S0_pff = ~((plm_out_acc_rmff==2'b10));
  assign plm_out_cns_d_shi1 = plm_out_cns_d_nsoftmax_compute_kernel_inst;
  assign plm_out_cns_radr_shi1 = plm_out_cns_radr_nsoftmax_store_output_inst;
  assign plm_out_cns_wadr_shi1 = plm_out_cns_wadr_nsoftmax_compute_kernel_inst;
  assign plm_out_cns_we_shi1 = plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_pff
      & plm_out_cns_S0_pff & plm_out_xor_rmff;
  assign plm_out_cns_S1 = (plm_out_acc_1_rmff!=2'b00);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cns_we_nsoftmax_compute_kernel_inst_buy <= 1'b0;
      plm_out_cns_ppidx <= 1'b0;
      plm_out_cns_ppown <= 2'b00;
      plm_out_cns_ppidx_1 <= 1'b0;
      plm_out_cns_ppown_1 <= 2'b00;
    end
    else begin
      plm_out_cns_we_nsoftmax_compute_kernel_inst_buy <= plm_out_cns_we_nsoftmax_compute_kernel_inst;
      plm_out_cns_ppidx <= plm_out_xor_rmff;
      plm_out_cns_ppown <= plm_out_acc_rmff;
      plm_out_cns_ppidx_1 <= plm_out_cns_ppidx_1 ^ plm_out_cns_PC1;
      plm_out_cns_ppown_1 <= plm_out_acc_1_rmff;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_plm_in_cns_bctl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_plm_in_cns_bctl (
  clk, rst, plm_in_cns_wadr_nsoftmax_load_input_inst, plm_in_cns_d_nsoftmax_load_input_inst,
      plm_in_cns_we_nsoftmax_load_input_inst, plm_in_cns_req_vz_nsoftmax_load_input_inst,
      plm_in_cns_radr_nsoftmax_compute_kernel_inst, plm_in_cns_q_nsoftmax_compute_kernel_inst,
      plm_in_cns_req_vz_nsoftmax_compute_kernel_inst, plm_out_cns_we_nsoftmax_compute_kernel_inst_buz,
      plm_in_cns_rls_lz_nsoftmax_load_input_inst_bud, plm_in_cns_rls_lz_nsoftmax_compute_kernel_inst_bud,
      plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud, plm_out_cns_rls_lz_nsoftmax_compute_kernel_inst_bud,
      plm_in_cns_S0, plm_in_cns_R0, plm_in_cns_S1, plm_in_cns_R1, plm_in_cns_d_shi0,
      plm_in_cns_d_shi1, plm_in_cns_q_sho0, plm_in_cns_q_sho1, plm_in_cns_radr_shi0,
      plm_in_cns_radr_shi1, plm_in_cns_wadr_shi0, plm_in_cns_wadr_shi1, plm_in_cns_we_shi0,
      plm_in_cns_we_shi1, plm_in_cns_S0_pff, plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_pff,
      plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud_pff
);
  input clk;
  input rst;
  input [6:0] plm_in_cns_wadr_nsoftmax_load_input_inst;
  input [31:0] plm_in_cns_d_nsoftmax_load_input_inst;
  input plm_in_cns_we_nsoftmax_load_input_inst;
  output plm_in_cns_req_vz_nsoftmax_load_input_inst;
  input [6:0] plm_in_cns_radr_nsoftmax_compute_kernel_inst;
  output [31:0] plm_in_cns_q_nsoftmax_compute_kernel_inst;
  output plm_in_cns_req_vz_nsoftmax_compute_kernel_inst;
  output plm_out_cns_we_nsoftmax_compute_kernel_inst_buz;
  input plm_in_cns_rls_lz_nsoftmax_load_input_inst_bud;
  input plm_in_cns_rls_lz_nsoftmax_compute_kernel_inst_bud;
  input plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud;
  input plm_out_cns_rls_lz_nsoftmax_compute_kernel_inst_bud;
  output plm_in_cns_S0;
  input plm_in_cns_R0;
  output plm_in_cns_S1;
  input plm_in_cns_R1;
  output [31:0] plm_in_cns_d_shi0;
  output [31:0] plm_in_cns_d_shi1;
  input [31:0] plm_in_cns_q_sho0;
  input [31:0] plm_in_cns_q_sho1;
  output [6:0] plm_in_cns_radr_shi0;
  output [6:0] plm_in_cns_radr_shi1;
  output [6:0] plm_in_cns_wadr_shi0;
  output [6:0] plm_in_cns_wadr_shi1;
  output plm_in_cns_we_shi0;
  output plm_in_cns_we_shi1;
  output plm_in_cns_S0_pff;
  output plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_pff;
  input plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud_pff;


  // Interconnect Declarations
  wire plm_in_cns_PC0;
  reg plm_in_cns_ppidx;
  reg [1:0] plm_in_cns_ppown;
  wire plm_in_cns_PC1;
  reg plm_in_cns_ppidx_1;
  reg [1:0] plm_in_cns_ppown_1;
  wire [1:0] plm_in_acc_rmff;
  wire [3:0] nl_plm_in_acc_rmff;
  wire plm_in_xor_rmff;
  wire [1:0] plm_in_acc_1_rmff;
  wire [3:0] nl_plm_in_acc_1_rmff;


  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_req_vz_nsoftmax_load_input_inst = plm_in_cns_R0;
  assign plm_in_cns_req_vz_nsoftmax_compute_kernel_inst = plm_in_cns_R1;
  assign plm_in_xor_rmff = plm_in_cns_ppidx ^ plm_in_cns_PC0;
  assign nl_plm_in_acc_rmff = plm_in_cns_ppown + conv_u2u_1_2(plm_in_cns_PC0) + conv_s2u_1_2(plm_in_cns_PC1);
  assign plm_in_acc_rmff = nl_plm_in_acc_rmff[1:0];
  assign plm_in_cns_PC0 = plm_in_cns_S0 & plm_in_cns_rls_lz_nsoftmax_load_input_inst_bud;
  assign nl_plm_in_acc_1_rmff = plm_in_cns_ppown_1 + conv_u2u_1_2(plm_in_cns_PC1)
      + conv_s2u_1_2(plm_in_cns_PC0);
  assign plm_in_acc_1_rmff = nl_plm_in_acc_1_rmff[1:0];
  assign plm_in_cns_PC1 = ((plm_in_cns_ppown_1!=2'b00)) & plm_in_cns_rls_lz_nsoftmax_compute_kernel_inst_bud;
  assign plm_in_cns_q_nsoftmax_compute_kernel_inst = MUX_v_32_2_2(plm_in_cns_q_sho0,
      plm_in_cns_q_sho1, plm_in_cns_ppidx_1);
  assign plm_in_cns_d_shi0 = plm_in_cns_d_nsoftmax_load_input_inst;
  assign plm_in_cns_radr_shi0 = plm_in_cns_radr_nsoftmax_compute_kernel_inst;
  assign plm_in_cns_wadr_shi0 = plm_in_cns_wadr_nsoftmax_load_input_inst;
  assign plm_in_cns_we_shi0 = plm_in_cns_we_nsoftmax_load_input_inst & plm_in_cns_S0_pff
      & (~ plm_in_xor_rmff);
  assign plm_in_cns_S0 = ~((plm_in_cns_ppown==2'b10));
  assign plm_in_cns_S0_pff = ~((plm_in_acc_rmff==2'b10));
  assign plm_in_cns_d_shi1 = plm_in_cns_d_nsoftmax_load_input_inst;
  assign plm_in_cns_radr_shi1 = plm_in_cns_radr_nsoftmax_compute_kernel_inst;
  assign plm_in_cns_wadr_shi1 = plm_in_cns_wadr_nsoftmax_load_input_inst;
  assign plm_in_cns_we_shi1 = plm_in_cns_we_nsoftmax_load_input_inst & plm_in_cns_S0_pff
      & plm_in_xor_rmff;
  assign plm_out_cns_we_nsoftmax_compute_kernel_inst_buz = plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud;
  assign plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_pff = plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud_pff;
  assign plm_in_cns_S1 = (plm_in_acc_1_rmff!=2'b00);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cns_ppidx <= 1'b0;
      plm_in_cns_ppown <= 2'b00;
      plm_in_cns_ppidx_1 <= 1'b0;
      plm_in_cns_ppown_1 <= 2'b00;
    end
    else begin
      plm_in_cns_ppidx <= plm_in_xor_rmff;
      plm_in_cns_ppown <= plm_in_acc_rmff;
      plm_in_cns_ppidx_1 <= plm_in_cns_ppidx_1 ^ plm_in_cns_PC1;
      plm_in_cns_ppown_1 <= plm_in_acc_1_rmff;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2u_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_unreg_hier
// ------------------------------------------------------------------


module esp_acc_softmax_unreg_hier (
  in_0, out_0
);
  input in_0;
  output out_0;



  // Interconnect Declarations for Component Instantiations 
  assign out_0 = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_7_32_128_128_32_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_7_32_128_128_32_1_gen
    (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [6:0] radr;
  output [31:0] q_d;
  input [6:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_store_output_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_store_output_fsm (
  clk, rst, store_output_wen, fsm_output, WAIT_FOR_CONFIG_LOOP_C_0_tr0, STORE_BATCH_LOOP_C_0_tr0
);
  input clk;
  input rst;
  input store_output_wen;
  output [6:0] fsm_output;
  reg [6:0] fsm_output;
  input WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  input STORE_BATCH_LOOP_C_0_tr0;


  // FSM State Type Declaration for esp_acc_softmax_softmax_store_output_store_output_store_output_fsm_1
  parameter
    WAIT_FOR_CONFIG_LOOP_C_0 = 3'd0,
    STORE_BATCH_LOOP_C_0 = 3'd1,
    store_output_rlp_C_0 = 3'd2,
    store_output_rlp_C_1 = 3'd3,
    store_output_rlp_C_2 = 3'd4,
    store_output_rlp_C_3 = 3'd5,
    PROCESS_DONE_LOOP_C_0 = 3'd6;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_softmax_softmax_store_output_store_output_store_output_fsm_1
    case (state_var)
      STORE_BATCH_LOOP_C_0 : begin
        fsm_output = 7'b0000010;
        if ( STORE_BATCH_LOOP_C_0_tr0 ) begin
          state_var_NS = STORE_BATCH_LOOP_C_0;
        end
        else begin
          state_var_NS = store_output_rlp_C_0;
        end
      end
      store_output_rlp_C_0 : begin
        fsm_output = 7'b0000100;
        state_var_NS = store_output_rlp_C_1;
      end
      store_output_rlp_C_1 : begin
        fsm_output = 7'b0001000;
        state_var_NS = store_output_rlp_C_2;
      end
      store_output_rlp_C_2 : begin
        fsm_output = 7'b0010000;
        state_var_NS = store_output_rlp_C_3;
      end
      store_output_rlp_C_3 : begin
        fsm_output = 7'b0100000;
        state_var_NS = PROCESS_DONE_LOOP_C_0;
      end
      PROCESS_DONE_LOOP_C_0 : begin
        fsm_output = 7'b1000000;
        state_var_NS = PROCESS_DONE_LOOP_C_0;
      end
      // WAIT_FOR_CONFIG_LOOP_C_0
      default : begin
        fsm_output = 7'b0000001;
        if ( WAIT_FOR_CONFIG_LOOP_C_0_tr0 ) begin
          state_var_NS = WAIT_FOR_CONFIG_LOOP_C_0;
        end
        else begin
          state_var_NS = STORE_BATCH_LOOP_C_0;
        end
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= WAIT_FOR_CONFIG_LOOP_C_0;
    end
    else if ( store_output_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_staller
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_staller (
  clk, rst, store_output_wen, store_output_wten, output_ready_ack_mioi_wen_comp,
      dma_write_ctrl_Push_mioi_wen_comp, dma_write_chnl_Push_mioi_wen_comp, plm_out_cns_req_obj_wen_comp
);
  input clk;
  input rst;
  output store_output_wen;
  output store_output_wten;
  input output_ready_ack_mioi_wen_comp;
  input dma_write_ctrl_Push_mioi_wen_comp;
  input dma_write_chnl_Push_mioi_wen_comp;
  input plm_out_cns_req_obj_wen_comp;


  // Interconnect Declarations
  reg store_output_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign store_output_wen = output_ready_ack_mioi_wen_comp & dma_write_ctrl_Push_mioi_wen_comp
      & dma_write_chnl_Push_mioi_wen_comp & plm_out_cns_req_obj_wen_comp;
  assign store_output_wten = store_output_wten_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      store_output_wten_reg <= 1'b0;
    end
    else begin
      store_output_wten_reg <= ~ store_output_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_req_obj_plm_out_cns_req_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_req_obj_plm_out_cns_req_wait_dp
    (
  clk, rst, plm_out_cns_req_obj_oswt, plm_out_cns_req_obj_wen_comp, plm_out_cns_req_obj_biwt,
      plm_out_cns_req_obj_bdwt, plm_out_cns_req_obj_bcwt
);
  input clk;
  input rst;
  input plm_out_cns_req_obj_oswt;
  output plm_out_cns_req_obj_wen_comp;
  input plm_out_cns_req_obj_biwt;
  input plm_out_cns_req_obj_bdwt;
  output plm_out_cns_req_obj_bcwt;
  reg plm_out_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_req_obj_wen_comp = (~ plm_out_cns_req_obj_oswt) | plm_out_cns_req_obj_biwt
      | plm_out_cns_req_obj_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cns_req_obj_bcwt <= 1'b0;
    end
    else begin
      plm_out_cns_req_obj_bcwt <= ~((~(plm_out_cns_req_obj_bcwt | plm_out_cns_req_obj_biwt))
          | plm_out_cns_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl
    (
  store_output_wen, plm_out_cns_req_obj_oswt, plm_out_cns_req_obj_vd, plm_out_cns_req_obj_biwt,
      plm_out_cns_req_obj_bdwt, plm_out_cns_req_obj_bcwt
);
  input store_output_wen;
  input plm_out_cns_req_obj_oswt;
  input plm_out_cns_req_obj_vd;
  output plm_out_cns_req_obj_biwt;
  output plm_out_cns_req_obj_bdwt;
  input plm_out_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_req_obj_bdwt = plm_out_cns_req_obj_oswt & store_output_wen;
  assign plm_out_cns_req_obj_biwt = plm_out_cns_req_obj_oswt & (~ plm_out_cns_req_obj_bcwt)
      & plm_out_cns_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl
    (
  store_output_wten, plm_out_cns_rls_obj_iswt0, plm_out_cns_rls_obj_ld_store_output_sct
);
  input store_output_wten;
  input plm_out_cns_rls_obj_iswt0;
  output plm_out_cns_rls_obj_ld_store_output_sct;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_rls_obj_ld_store_output_sct = plm_out_cns_rls_obj_iswt0 & (~
      store_output_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_1_plm_out_cns_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_1_plm_out_cns_wait_dp
    (
  clk, rst, plm_out_cnsi_q_d, plm_out_cnsi_q_d_mxwt, plm_out_cnsi_biwt, plm_out_cnsi_bdwt
);
  input clk;
  input rst;
  input [31:0] plm_out_cnsi_q_d;
  output [31:0] plm_out_cnsi_q_d_mxwt;
  input plm_out_cnsi_biwt;
  input plm_out_cnsi_bdwt;


  // Interconnect Declarations
  reg plm_out_cnsi_bcwt;
  reg [31:0] plm_out_cnsi_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cnsi_q_d_mxwt = MUX_v_32_2_2(plm_out_cnsi_q_d, plm_out_cnsi_q_d_bfwt,
      plm_out_cnsi_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cnsi_bcwt <= 1'b0;
    end
    else begin
      plm_out_cnsi_bcwt <= ~((~(plm_out_cnsi_bcwt | plm_out_cnsi_biwt)) | plm_out_cnsi_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( plm_out_cnsi_biwt ) begin
      plm_out_cnsi_q_d_bfwt <= plm_out_cnsi_q_d;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_1_plm_out_cns_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_1_plm_out_cns_wait_ctrl
    (
  store_output_wen, store_output_wten, plm_out_cnsi_oswt, plm_out_cnsi_biwt, plm_out_cnsi_bdwt,
      plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_store_output_sct, plm_out_cnsi_oswt_pff
);
  input store_output_wen;
  input store_output_wten;
  input plm_out_cnsi_oswt;
  output plm_out_cnsi_biwt;
  output plm_out_cnsi_bdwt;
  output plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_store_output_sct;
  input plm_out_cnsi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cnsi_bdwt = plm_out_cnsi_oswt & store_output_wen;
  assign plm_out_cnsi_biwt = (~ store_output_wten) & plm_out_cnsi_oswt;
  assign plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_store_output_sct = plm_out_cnsi_oswt_pff
      & store_output_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp
    (
  clk, rst, dma_write_chnl_Push_mioi_oswt, dma_write_chnl_Push_mioi_wen_comp, dma_write_chnl_Push_mioi_m_rsc_dat_store_output,
      dma_write_chnl_Push_mioi_m_rsc_dat, dma_write_chnl_Push_mioi_biwt, dma_write_chnl_Push_mioi_bdwt,
      dma_write_chnl_Push_mioi_bcwt, dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
);
  input clk;
  input rst;
  input dma_write_chnl_Push_mioi_oswt;
  output dma_write_chnl_Push_mioi_wen_comp;
  input [63:0] dma_write_chnl_Push_mioi_m_rsc_dat_store_output;
  output [63:0] dma_write_chnl_Push_mioi_m_rsc_dat;
  input dma_write_chnl_Push_mioi_biwt;
  input dma_write_chnl_Push_mioi_bdwt;
  output dma_write_chnl_Push_mioi_bcwt;
  reg dma_write_chnl_Push_mioi_bcwt;
  input dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dma_write_chnl_Push_mioi_wen_comp = (~ dma_write_chnl_Push_mioi_oswt) |
      dma_write_chnl_Push_mioi_biwt | dma_write_chnl_Push_mioi_bcwt;
  assign dma_write_chnl_Push_mioi_m_rsc_dat = {dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff)
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff) , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff) , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff) , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff)
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff) , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff) , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff) , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , (dma_write_chnl_Push_mioi_m_rsc_dat_store_output[31:0])};
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_chnl_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_write_chnl_Push_mioi_bcwt <= ~((~(dma_write_chnl_Push_mioi_bcwt | dma_write_chnl_Push_mioi_biwt))
          | dma_write_chnl_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl
    (
  store_output_wen, dma_write_chnl_Push_mioi_oswt, dma_write_chnl_Push_mioi_biwt,
      dma_write_chnl_Push_mioi_bdwt, dma_write_chnl_Push_mioi_bcwt, dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld,
      dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff, dma_write_chnl_Push_mioi_oswt_pff
);
  input store_output_wen;
  input dma_write_chnl_Push_mioi_oswt;
  output dma_write_chnl_Push_mioi_biwt;
  output dma_write_chnl_Push_mioi_bdwt;
  input dma_write_chnl_Push_mioi_bcwt;
  input dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld;
  output dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff;
  input dma_write_chnl_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dma_write_chnl_Push_mioi_bdwt = dma_write_chnl_Push_mioi_oswt & store_output_wen;
  assign dma_write_chnl_Push_mioi_biwt = dma_write_chnl_Push_mioi_oswt & (~ dma_write_chnl_Push_mioi_bcwt)
      & dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld;
  assign dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff = dma_write_chnl_Push_mioi_oswt_pff
      & store_output_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp
    (
  clk, rst, dma_write_ctrl_Push_mioi_oswt, dma_write_ctrl_Push_mioi_wen_comp, dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output,
      dma_write_ctrl_Push_mioi_m_index_rsc_dat, dma_write_ctrl_Push_mioi_biwt, dma_write_ctrl_Push_mioi_bdwt,
      dma_write_ctrl_Push_mioi_bcwt, dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_pff
);
  input clk;
  input rst;
  input dma_write_ctrl_Push_mioi_oswt;
  output dma_write_ctrl_Push_mioi_wen_comp;
  input [31:0] dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output;
  output [31:0] dma_write_ctrl_Push_mioi_m_index_rsc_dat;
  input dma_write_ctrl_Push_mioi_biwt;
  input dma_write_ctrl_Push_mioi_bdwt;
  output dma_write_ctrl_Push_mioi_bcwt;
  reg dma_write_ctrl_Push_mioi_bcwt;
  input dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dma_write_ctrl_Push_mioi_wen_comp = (~ dma_write_ctrl_Push_mioi_oswt) |
      dma_write_ctrl_Push_mioi_biwt | dma_write_ctrl_Push_mioi_bcwt;
  assign dma_write_ctrl_Push_mioi_m_index_rsc_dat = {(dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output[31:7])
      , (~ dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_pff) , (~ dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_pff)
      , (~ dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_pff) , (~ dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_pff)
      , (~ dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_pff) , (~ dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_pff)
      , (~ dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_pff)};
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_ctrl_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_write_ctrl_Push_mioi_bcwt <= ~((~(dma_write_ctrl_Push_mioi_bcwt | dma_write_ctrl_Push_mioi_biwt))
          | dma_write_ctrl_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl
    (
  store_output_wen, dma_write_ctrl_Push_mioi_oswt, dma_write_ctrl_Push_mioi_biwt,
      dma_write_ctrl_Push_mioi_bdwt, dma_write_ctrl_Push_mioi_bcwt, dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld,
      dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_pff, dma_write_ctrl_Push_mioi_oswt_pff
);
  input store_output_wen;
  input dma_write_ctrl_Push_mioi_oswt;
  output dma_write_ctrl_Push_mioi_biwt;
  output dma_write_ctrl_Push_mioi_bdwt;
  input dma_write_ctrl_Push_mioi_bcwt;
  input dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  output dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_pff;
  input dma_write_ctrl_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dma_write_ctrl_Push_mioi_bdwt = dma_write_ctrl_Push_mioi_oswt & store_output_wen;
  assign dma_write_ctrl_Push_mioi_biwt = dma_write_ctrl_Push_mioi_oswt & (~ dma_write_ctrl_Push_mioi_bcwt)
      & dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  assign dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_pff = dma_write_ctrl_Push_mioi_oswt_pff
      & store_output_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_output_ready_ack_mioi_output_ready_ack_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_output_ready_ack_mioi_output_ready_ack_mio_wait_dp
    (
  clk, rst, output_ready_ack_mioi_oswt, output_ready_ack_mioi_wen_comp, output_ready_ack_mioi_biwt,
      output_ready_ack_mioi_bdwt, output_ready_ack_mioi_bcwt
);
  input clk;
  input rst;
  input output_ready_ack_mioi_oswt;
  output output_ready_ack_mioi_wen_comp;
  input output_ready_ack_mioi_biwt;
  input output_ready_ack_mioi_bdwt;
  output output_ready_ack_mioi_bcwt;
  reg output_ready_ack_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign output_ready_ack_mioi_wen_comp = (~ output_ready_ack_mioi_oswt) | output_ready_ack_mioi_biwt
      | output_ready_ack_mioi_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      output_ready_ack_mioi_bcwt <= 1'b0;
    end
    else begin
      output_ready_ack_mioi_bcwt <= ~((~(output_ready_ack_mioi_bcwt | output_ready_ack_mioi_biwt))
          | output_ready_ack_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_output_ready_ack_mioi_output_ready_ack_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_output_ready_ack_mioi_output_ready_ack_mio_wait_ctrl
    (
  store_output_wen, output_ready_ack_mioi_oswt, output_ready_ack_mioi_biwt, output_ready_ack_mioi_bdwt,
      output_ready_ack_mioi_bcwt, output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_output_sct,
      output_ready_ack_mioi_ccs_ccore_done_sync_vld, output_ready_ack_mioi_oswt_pff
);
  input store_output_wen;
  input output_ready_ack_mioi_oswt;
  output output_ready_ack_mioi_biwt;
  output output_ready_ack_mioi_bdwt;
  input output_ready_ack_mioi_bcwt;
  output output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_output_sct;
  input output_ready_ack_mioi_ccs_ccore_done_sync_vld;
  input output_ready_ack_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign output_ready_ack_mioi_bdwt = output_ready_ack_mioi_oswt & store_output_wen;
  assign output_ready_ack_mioi_biwt = output_ready_ack_mioi_oswt & (~ output_ready_ack_mioi_bcwt)
      & output_ready_ack_mioi_ccs_ccore_done_sync_vld;
  assign output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_output_sct = output_ready_ack_mioi_oswt_pff
      & store_output_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_35_7_32_128_128_32_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_35_7_32_128_128_32_1_gen
    (
  we, d, wadr, d_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [31:0] d;
  output [6:0] wadr;
  input [31:0] d_d;
  input [6:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_7_32_128_128_32_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_7_32_128_128_32_1_gen
    (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [31:0] q;
  output [6:0] radr;
  output [31:0] q_d;
  input [6:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_17_7_67_128_128_67_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_17_7_67_128_128_67_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [66:0] q;
  output [6:0] radr;
  output we;
  output [66:0] d;
  output [6:0] wadr;
  input clken_d;
  input [66:0] d_d;
  output [66:0] q_d;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_compute_kernel_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_compute_kernel_fsm (
  clk, rst, compute_kernel_wen, fsm_output, WAIT_FOR_CONFIG_LOOP_C_0_tr0, COMPUTE_BATCH_LOOP_C_0_tr0
);
  input clk;
  input rst;
  input compute_kernel_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;
  input WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  input COMPUTE_BATCH_LOOP_C_0_tr0;


  // FSM State Type Declaration for esp_acc_softmax_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_1
  parameter
    WAIT_FOR_CONFIG_LOOP_C_0 = 2'd0,
    COMPUTE_BATCH_LOOP_C_0 = 2'd1,
    PROCESS_DONE_LOOP_C_0 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_softmax_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_1
    case (state_var)
      COMPUTE_BATCH_LOOP_C_0 : begin
        fsm_output = 3'b010;
        if ( COMPUTE_BATCH_LOOP_C_0_tr0 ) begin
          state_var_NS = COMPUTE_BATCH_LOOP_C_0;
        end
        else begin
          state_var_NS = PROCESS_DONE_LOOP_C_0;
        end
      end
      PROCESS_DONE_LOOP_C_0 : begin
        fsm_output = 3'b100;
        state_var_NS = PROCESS_DONE_LOOP_C_0;
      end
      // WAIT_FOR_CONFIG_LOOP_C_0
      default : begin
        fsm_output = 3'b001;
        if ( WAIT_FOR_CONFIG_LOOP_C_0_tr0 ) begin
          state_var_NS = WAIT_FOR_CONFIG_LOOP_C_0;
        end
        else begin
          state_var_NS = COMPUTE_BATCH_LOOP_C_0;
        end
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= WAIT_FOR_CONFIG_LOOP_C_0;
    end
    else if ( compute_kernel_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_staller
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_staller (
  clk, rst, compute_kernel_wen, compute_kernel_wten, input_ready_ack_mioi_wen_comp,
      output_ready_req_mioi_wen_comp, plm_in_cns_req_obj_wen_comp, plm_out_cns_req_obj_wen_comp
);
  input clk;
  input rst;
  output compute_kernel_wen;
  output compute_kernel_wten;
  input input_ready_ack_mioi_wen_comp;
  input output_ready_req_mioi_wen_comp;
  input plm_in_cns_req_obj_wen_comp;
  input plm_out_cns_req_obj_wen_comp;


  // Interconnect Declarations
  reg compute_kernel_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign compute_kernel_wen = input_ready_ack_mioi_wen_comp & output_ready_req_mioi_wen_comp
      & plm_in_cns_req_obj_wen_comp & plm_out_cns_req_obj_wen_comp;
  assign compute_kernel_wten = compute_kernel_wten_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      compute_kernel_wten_reg <= 1'b0;
    end
    else begin
      compute_kernel_wten_reg <= ~ compute_kernel_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_req_obj_plm_out_cns_req_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_req_obj_plm_out_cns_req_wait_dp
    (
  clk, rst, plm_out_cns_req_obj_oswt, plm_out_cns_req_obj_wen_comp, plm_out_cns_req_obj_biwt,
      plm_out_cns_req_obj_bdwt, plm_out_cns_req_obj_bcwt
);
  input clk;
  input rst;
  input plm_out_cns_req_obj_oswt;
  output plm_out_cns_req_obj_wen_comp;
  input plm_out_cns_req_obj_biwt;
  input plm_out_cns_req_obj_bdwt;
  output plm_out_cns_req_obj_bcwt;
  reg plm_out_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_req_obj_wen_comp = (~ plm_out_cns_req_obj_oswt) | plm_out_cns_req_obj_biwt
      | plm_out_cns_req_obj_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cns_req_obj_bcwt <= 1'b0;
    end
    else begin
      plm_out_cns_req_obj_bcwt <= ~((~(plm_out_cns_req_obj_bcwt | plm_out_cns_req_obj_biwt))
          | plm_out_cns_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl
    (
  compute_kernel_wen, plm_out_cns_req_obj_oswt, plm_out_cns_req_obj_vd, plm_out_cns_req_obj_biwt,
      plm_out_cns_req_obj_bdwt, plm_out_cns_req_obj_bcwt
);
  input compute_kernel_wen;
  input plm_out_cns_req_obj_oswt;
  input plm_out_cns_req_obj_vd;
  output plm_out_cns_req_obj_biwt;
  output plm_out_cns_req_obj_bdwt;
  input plm_out_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_req_obj_bdwt = plm_out_cns_req_obj_oswt & compute_kernel_wen;
  assign plm_out_cns_req_obj_biwt = plm_out_cns_req_obj_oswt & (~ plm_out_cns_req_obj_bcwt)
      & plm_out_cns_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_req_obj_plm_in_cns_req_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_req_obj_plm_in_cns_req_wait_dp
    (
  clk, rst, plm_in_cns_req_obj_oswt, plm_in_cns_req_obj_wen_comp, plm_in_cns_req_obj_biwt,
      plm_in_cns_req_obj_bdwt, plm_in_cns_req_obj_bcwt
);
  input clk;
  input rst;
  input plm_in_cns_req_obj_oswt;
  output plm_in_cns_req_obj_wen_comp;
  input plm_in_cns_req_obj_biwt;
  input plm_in_cns_req_obj_bdwt;
  output plm_in_cns_req_obj_bcwt;
  reg plm_in_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_req_obj_wen_comp = (~ plm_in_cns_req_obj_oswt) | plm_in_cns_req_obj_biwt
      | plm_in_cns_req_obj_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cns_req_obj_bcwt <= 1'b0;
    end
    else begin
      plm_in_cns_req_obj_bcwt <= ~((~(plm_in_cns_req_obj_bcwt | plm_in_cns_req_obj_biwt))
          | plm_in_cns_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl
    (
  compute_kernel_wen, plm_in_cns_req_obj_oswt, plm_in_cns_req_obj_vd, plm_in_cns_req_obj_biwt,
      plm_in_cns_req_obj_bdwt, plm_in_cns_req_obj_bcwt
);
  input compute_kernel_wen;
  input plm_in_cns_req_obj_oswt;
  input plm_in_cns_req_obj_vd;
  output plm_in_cns_req_obj_biwt;
  output plm_in_cns_req_obj_bdwt;
  input plm_in_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_req_obj_bdwt = plm_in_cns_req_obj_oswt & compute_kernel_wen;
  assign plm_in_cns_req_obj_biwt = plm_in_cns_req_obj_oswt & (~ plm_in_cns_req_obj_bcwt)
      & plm_in_cns_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl
    (
  compute_kernel_wten, plm_in_cns_rls_obj_iswt0, plm_in_cns_rls_obj_ld_compute_kernel_sct
);
  input compute_kernel_wten;
  input plm_in_cns_rls_obj_iswt0;
  output plm_in_cns_rls_obj_ld_compute_kernel_sct;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_rls_obj_ld_compute_kernel_sct = plm_in_cns_rls_obj_iswt0 & (~
      compute_kernel_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl
    (
  compute_kernel_wten, plm_out_cns_rls_obj_iswt0, plm_out_cns_rls_obj_ld_compute_kernel_sct
);
  input compute_kernel_wten;
  input plm_out_cns_rls_obj_iswt0;
  output plm_out_cns_rls_obj_ld_compute_kernel_sct;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cns_rls_obj_ld_compute_kernel_sct = plm_out_cns_rls_obj_iswt0 &
      (~ compute_kernel_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi_1_plm_out_cns_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi_1_plm_out_cns_wait_ctrl
    (
  plm_out_cnsi_we_d_compute_kernel_sct_pff, plm_out_cnsi_iswt0_pff, compute_kernel_wten_pff
);
  output plm_out_cnsi_we_d_compute_kernel_sct_pff;
  input plm_out_cnsi_iswt0_pff;
  input compute_kernel_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cnsi_we_d_compute_kernel_sct_pff = plm_out_cnsi_iswt0_pff & (~ compute_kernel_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_1_plm_in_cns_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_1_plm_in_cns_wait_dp
    (
  clk, rst, plm_in_cnsi_q_d, plm_in_cnsi_q_d_mxwt, plm_in_cnsi_biwt, plm_in_cnsi_bdwt
);
  input clk;
  input rst;
  input [31:0] plm_in_cnsi_q_d;
  output [31:0] plm_in_cnsi_q_d_mxwt;
  input plm_in_cnsi_biwt;
  input plm_in_cnsi_bdwt;


  // Interconnect Declarations
  reg plm_in_cnsi_bcwt;
  reg [31:0] plm_in_cnsi_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cnsi_q_d_mxwt = MUX_v_32_2_2(plm_in_cnsi_q_d, plm_in_cnsi_q_d_bfwt,
      plm_in_cnsi_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cnsi_bcwt <= 1'b0;
    end
    else begin
      plm_in_cnsi_bcwt <= ~((~(plm_in_cnsi_bcwt | plm_in_cnsi_biwt)) | plm_in_cnsi_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( plm_in_cnsi_biwt ) begin
      plm_in_cnsi_q_d_bfwt <= plm_in_cnsi_q_d;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_1_plm_in_cns_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_1_plm_in_cns_wait_ctrl
    (
  compute_kernel_wen, compute_kernel_wten, plm_in_cnsi_oswt, plm_in_cnsi_biwt, plm_in_cnsi_bdwt,
      plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_compute_kernel_sct, plm_in_cnsi_oswt_pff
);
  input compute_kernel_wen;
  input compute_kernel_wten;
  input plm_in_cnsi_oswt;
  output plm_in_cnsi_biwt;
  output plm_in_cnsi_bdwt;
  output plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_compute_kernel_sct;
  input plm_in_cnsi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cnsi_bdwt = plm_in_cnsi_oswt & compute_kernel_wen;
  assign plm_in_cnsi_biwt = (~ compute_kernel_wten) & plm_in_cnsi_oswt;
  assign plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_compute_kernel_sct = plm_in_cnsi_oswt_pff
      & compute_kernel_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_req_mioi_output_ready_req_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_req_mioi_output_ready_req_mio_wait_dp
    (
  clk, rst, output_ready_req_mioi_oswt, output_ready_req_mioi_wen_comp, output_ready_req_mioi_biwt,
      output_ready_req_mioi_bdwt, output_ready_req_mioi_bcwt
);
  input clk;
  input rst;
  input output_ready_req_mioi_oswt;
  output output_ready_req_mioi_wen_comp;
  input output_ready_req_mioi_biwt;
  input output_ready_req_mioi_bdwt;
  output output_ready_req_mioi_bcwt;
  reg output_ready_req_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign output_ready_req_mioi_wen_comp = (~ output_ready_req_mioi_oswt) | output_ready_req_mioi_biwt
      | output_ready_req_mioi_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      output_ready_req_mioi_bcwt <= 1'b0;
    end
    else begin
      output_ready_req_mioi_bcwt <= ~((~(output_ready_req_mioi_bcwt | output_ready_req_mioi_biwt))
          | output_ready_req_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_req_mioi_output_ready_req_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_req_mioi_output_ready_req_mio_wait_ctrl
    (
  compute_kernel_wen, output_ready_req_mioi_oswt, output_ready_req_mioi_biwt, output_ready_req_mioi_bdwt,
      output_ready_req_mioi_bcwt, output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct,
      output_ready_req_mioi_ccs_ccore_done_sync_vld, output_ready_req_mioi_oswt_pff
);
  input compute_kernel_wen;
  input output_ready_req_mioi_oswt;
  output output_ready_req_mioi_biwt;
  output output_ready_req_mioi_bdwt;
  input output_ready_req_mioi_bcwt;
  output output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct;
  input output_ready_req_mioi_ccs_ccore_done_sync_vld;
  input output_ready_req_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign output_ready_req_mioi_bdwt = output_ready_req_mioi_oswt & compute_kernel_wen;
  assign output_ready_req_mioi_biwt = output_ready_req_mioi_oswt & (~ output_ready_req_mioi_bcwt)
      & output_ready_req_mioi_ccs_ccore_done_sync_vld;
  assign output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct = output_ready_req_mioi_oswt_pff
      & compute_kernel_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_ack_mioi_input_ready_ack_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_ack_mioi_input_ready_ack_mio_wait_dp
    (
  clk, rst, input_ready_ack_mioi_oswt, input_ready_ack_mioi_wen_comp, input_ready_ack_mioi_biwt,
      input_ready_ack_mioi_bdwt, input_ready_ack_mioi_bcwt
);
  input clk;
  input rst;
  input input_ready_ack_mioi_oswt;
  output input_ready_ack_mioi_wen_comp;
  input input_ready_ack_mioi_biwt;
  input input_ready_ack_mioi_bdwt;
  output input_ready_ack_mioi_bcwt;
  reg input_ready_ack_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign input_ready_ack_mioi_wen_comp = (~ input_ready_ack_mioi_oswt) | input_ready_ack_mioi_biwt
      | input_ready_ack_mioi_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      input_ready_ack_mioi_bcwt <= 1'b0;
    end
    else begin
      input_ready_ack_mioi_bcwt <= ~((~(input_ready_ack_mioi_bcwt | input_ready_ack_mioi_biwt))
          | input_ready_ack_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_ack_mioi_input_ready_ack_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_ack_mioi_input_ready_ack_mio_wait_ctrl
    (
  compute_kernel_wen, input_ready_ack_mioi_oswt, input_ready_ack_mioi_biwt, input_ready_ack_mioi_bdwt,
      input_ready_ack_mioi_bcwt, input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct,
      input_ready_ack_mioi_ccs_ccore_done_sync_vld, input_ready_ack_mioi_oswt_pff
);
  input compute_kernel_wen;
  input input_ready_ack_mioi_oswt;
  output input_ready_ack_mioi_biwt;
  output input_ready_ack_mioi_bdwt;
  input input_ready_ack_mioi_bcwt;
  output input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct;
  input input_ready_ack_mioi_ccs_ccore_done_sync_vld;
  input input_ready_ack_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign input_ready_ack_mioi_bdwt = input_ready_ack_mioi_oswt & compute_kernel_wen;
  assign input_ready_ack_mioi_biwt = input_ready_ack_mioi_oswt & (~ input_ready_ack_mioi_bcwt)
      & input_ready_ack_mioi_ccs_ccore_done_sync_vld;
  assign input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct = input_ready_ack_mioi_oswt_pff
      & compute_kernel_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_33_7_32_128_128_32_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_33_7_32_128_128_32_1_gen
    (
  we, d, wadr, d_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [31:0] d;
  output [6:0] wadr;
  input [31:0] d_d;
  input [6:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_load_input_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_load_input_fsm (
  clk, rst, load_input_wen, fsm_output, WAIT_FOR_CONFIG_LOOP_C_0_tr0, LOAD_BATCH_LOOP_C_0_tr0
);
  input clk;
  input rst;
  input load_input_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;
  input WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  input LOAD_BATCH_LOOP_C_0_tr0;


  // FSM State Type Declaration for esp_acc_softmax_softmax_load_input_load_input_load_input_fsm_1
  parameter
    WAIT_FOR_CONFIG_LOOP_C_0 = 2'd0,
    LOAD_BATCH_LOOP_C_0 = 2'd1,
    PROCESS_DONE_LOOP_C_0 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_softmax_softmax_load_input_load_input_load_input_fsm_1
    case (state_var)
      LOAD_BATCH_LOOP_C_0 : begin
        fsm_output = 3'b010;
        if ( LOAD_BATCH_LOOP_C_0_tr0 ) begin
          state_var_NS = LOAD_BATCH_LOOP_C_0;
        end
        else begin
          state_var_NS = PROCESS_DONE_LOOP_C_0;
        end
      end
      PROCESS_DONE_LOOP_C_0 : begin
        fsm_output = 3'b100;
        state_var_NS = PROCESS_DONE_LOOP_C_0;
      end
      // WAIT_FOR_CONFIG_LOOP_C_0
      default : begin
        fsm_output = 3'b001;
        if ( WAIT_FOR_CONFIG_LOOP_C_0_tr0 ) begin
          state_var_NS = WAIT_FOR_CONFIG_LOOP_C_0;
        end
        else begin
          state_var_NS = LOAD_BATCH_LOOP_C_0;
        end
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= WAIT_FOR_CONFIG_LOOP_C_0;
    end
    else if ( load_input_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_staller
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_staller (
  clk, rst, load_input_wen, load_input_wten, dma_read_ctrl_Push_mioi_wen_comp, dma_read_chnl_Pop_mioi_wen_comp,
      input_ready_req_mioi_wen_comp, plm_in_cns_req_obj_wen_comp
);
  input clk;
  input rst;
  output load_input_wen;
  output load_input_wten;
  input dma_read_ctrl_Push_mioi_wen_comp;
  input dma_read_chnl_Pop_mioi_wen_comp;
  input input_ready_req_mioi_wen_comp;
  input plm_in_cns_req_obj_wen_comp;


  // Interconnect Declarations
  reg load_input_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign load_input_wen = dma_read_ctrl_Push_mioi_wen_comp & dma_read_chnl_Pop_mioi_wen_comp
      & input_ready_req_mioi_wen_comp & plm_in_cns_req_obj_wen_comp;
  assign load_input_wten = load_input_wten_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      load_input_wten_reg <= 1'b0;
    end
    else begin
      load_input_wten_reg <= ~ load_input_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_req_obj_plm_in_cns_req_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_req_obj_plm_in_cns_req_wait_dp
    (
  clk, rst, plm_in_cns_req_obj_oswt, plm_in_cns_req_obj_wen_comp, plm_in_cns_req_obj_biwt,
      plm_in_cns_req_obj_bdwt, plm_in_cns_req_obj_bcwt
);
  input clk;
  input rst;
  input plm_in_cns_req_obj_oswt;
  output plm_in_cns_req_obj_wen_comp;
  input plm_in_cns_req_obj_biwt;
  input plm_in_cns_req_obj_bdwt;
  output plm_in_cns_req_obj_bcwt;
  reg plm_in_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_req_obj_wen_comp = (~ plm_in_cns_req_obj_oswt) | plm_in_cns_req_obj_biwt
      | plm_in_cns_req_obj_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cns_req_obj_bcwt <= 1'b0;
    end
    else begin
      plm_in_cns_req_obj_bcwt <= ~((~(plm_in_cns_req_obj_bcwt | plm_in_cns_req_obj_biwt))
          | plm_in_cns_req_obj_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl
    (
  load_input_wen, plm_in_cns_req_obj_oswt, plm_in_cns_req_obj_vd, plm_in_cns_req_obj_biwt,
      plm_in_cns_req_obj_bdwt, plm_in_cns_req_obj_bcwt
);
  input load_input_wen;
  input plm_in_cns_req_obj_oswt;
  input plm_in_cns_req_obj_vd;
  output plm_in_cns_req_obj_biwt;
  output plm_in_cns_req_obj_bdwt;
  input plm_in_cns_req_obj_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_req_obj_bdwt = plm_in_cns_req_obj_oswt & load_input_wen;
  assign plm_in_cns_req_obj_biwt = plm_in_cns_req_obj_oswt & (~ plm_in_cns_req_obj_bcwt)
      & plm_in_cns_req_obj_vd;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl
    (
  load_input_wten, plm_in_cns_rls_obj_iswt0, plm_in_cns_rls_obj_ld_load_input_sct
);
  input load_input_wten;
  input plm_in_cns_rls_obj_iswt0;
  output plm_in_cns_rls_obj_ld_load_input_sct;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cns_rls_obj_ld_load_input_sct = plm_in_cns_rls_obj_iswt0 & (~ load_input_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi_1_plm_in_cns_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi_1_plm_in_cns_wait_ctrl
    (
  plm_in_cnsi_we_d_load_input_sct_pff, plm_in_cnsi_iswt0_pff, load_input_wten_pff
);
  output plm_in_cnsi_we_d_load_input_sct_pff;
  input plm_in_cnsi_iswt0_pff;
  input load_input_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cnsi_we_d_load_input_sct_pff = plm_in_cnsi_iswt0_pff & (~ load_input_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_input_ready_req_mioi_input_ready_req_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_input_ready_req_mioi_input_ready_req_mio_wait_dp
    (
  clk, rst, input_ready_req_mioi_oswt, input_ready_req_mioi_wen_comp, input_ready_req_mioi_biwt,
      input_ready_req_mioi_bdwt, input_ready_req_mioi_bcwt
);
  input clk;
  input rst;
  input input_ready_req_mioi_oswt;
  output input_ready_req_mioi_wen_comp;
  input input_ready_req_mioi_biwt;
  input input_ready_req_mioi_bdwt;
  output input_ready_req_mioi_bcwt;
  reg input_ready_req_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign input_ready_req_mioi_wen_comp = (~ input_ready_req_mioi_oswt) | input_ready_req_mioi_biwt
      | input_ready_req_mioi_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      input_ready_req_mioi_bcwt <= 1'b0;
    end
    else begin
      input_ready_req_mioi_bcwt <= ~((~(input_ready_req_mioi_bcwt | input_ready_req_mioi_biwt))
          | input_ready_req_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_input_ready_req_mioi_input_ready_req_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_input_ready_req_mioi_input_ready_req_mio_wait_ctrl
    (
  load_input_wen, input_ready_req_mioi_oswt, input_ready_req_mioi_biwt, input_ready_req_mioi_bdwt,
      input_ready_req_mioi_bcwt, input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_input_sct,
      input_ready_req_mioi_ccs_ccore_done_sync_vld, input_ready_req_mioi_oswt_pff
);
  input load_input_wen;
  input input_ready_req_mioi_oswt;
  output input_ready_req_mioi_biwt;
  output input_ready_req_mioi_bdwt;
  input input_ready_req_mioi_bcwt;
  output input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_input_sct;
  input input_ready_req_mioi_ccs_ccore_done_sync_vld;
  input input_ready_req_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign input_ready_req_mioi_bdwt = input_ready_req_mioi_oswt & load_input_wen;
  assign input_ready_req_mioi_biwt = input_ready_req_mioi_oswt & (~ input_ready_req_mioi_bcwt)
      & input_ready_req_mioi_ccs_ccore_done_sync_vld;
  assign input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_input_sct = input_ready_req_mioi_oswt_pff
      & load_input_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp
    (
  clk, rst, dma_read_chnl_Pop_mioi_oswt, dma_read_chnl_Pop_mioi_wen_comp, dma_read_chnl_Pop_mioi_return_rsc_z_mxwt,
      dma_read_chnl_Pop_mioi_return_rsc_z, dma_read_chnl_Pop_mioi_biwt, dma_read_chnl_Pop_mioi_bdwt,
      dma_read_chnl_Pop_mioi_bcwt
);
  input clk;
  input rst;
  input dma_read_chnl_Pop_mioi_oswt;
  output dma_read_chnl_Pop_mioi_wen_comp;
  output [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt;
  input [63:0] dma_read_chnl_Pop_mioi_return_rsc_z;
  input dma_read_chnl_Pop_mioi_biwt;
  input dma_read_chnl_Pop_mioi_bdwt;
  output dma_read_chnl_Pop_mioi_bcwt;
  reg dma_read_chnl_Pop_mioi_bcwt;


  // Interconnect Declarations
  reg [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_bfwt_31_0;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_chnl_Pop_mioi_wen_comp = (~ dma_read_chnl_Pop_mioi_oswt) | dma_read_chnl_Pop_mioi_biwt
      | dma_read_chnl_Pop_mioi_bcwt;
  assign dma_read_chnl_Pop_mioi_return_rsc_z_mxwt = MUX_v_32_2_2((dma_read_chnl_Pop_mioi_return_rsc_z[31:0]),
      dma_read_chnl_Pop_mioi_return_rsc_z_bfwt_31_0, dma_read_chnl_Pop_mioi_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_chnl_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_read_chnl_Pop_mioi_bcwt <= ~((~(dma_read_chnl_Pop_mioi_bcwt | dma_read_chnl_Pop_mioi_biwt))
          | dma_read_chnl_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( dma_read_chnl_Pop_mioi_biwt ) begin
      dma_read_chnl_Pop_mioi_return_rsc_z_bfwt_31_0 <= dma_read_chnl_Pop_mioi_return_rsc_z[31:0];
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl
    (
  load_input_wen, dma_read_chnl_Pop_mioi_oswt, dma_read_chnl_Pop_mioi_biwt, dma_read_chnl_Pop_mioi_bdwt,
      dma_read_chnl_Pop_mioi_bcwt, dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct,
      dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld, dma_read_chnl_Pop_mioi_oswt_pff
);
  input load_input_wen;
  input dma_read_chnl_Pop_mioi_oswt;
  output dma_read_chnl_Pop_mioi_biwt;
  output dma_read_chnl_Pop_mioi_bdwt;
  input dma_read_chnl_Pop_mioi_bcwt;
  output dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct;
  input dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld;
  input dma_read_chnl_Pop_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dma_read_chnl_Pop_mioi_bdwt = dma_read_chnl_Pop_mioi_oswt & load_input_wen;
  assign dma_read_chnl_Pop_mioi_biwt = dma_read_chnl_Pop_mioi_oswt & (~ dma_read_chnl_Pop_mioi_bcwt)
      & dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld;
  assign dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct = dma_read_chnl_Pop_mioi_oswt_pff
      & load_input_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp
    (
  clk, rst, dma_read_ctrl_Push_mioi_oswt, dma_read_ctrl_Push_mioi_wen_comp, dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input,
      dma_read_ctrl_Push_mioi_m_index_rsc_dat, dma_read_ctrl_Push_mioi_biwt, dma_read_ctrl_Push_mioi_bdwt,
      dma_read_ctrl_Push_mioi_bcwt, dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_pff
);
  input clk;
  input rst;
  input dma_read_ctrl_Push_mioi_oswt;
  output dma_read_ctrl_Push_mioi_wen_comp;
  input [31:0] dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input;
  output [31:0] dma_read_ctrl_Push_mioi_m_index_rsc_dat;
  input dma_read_ctrl_Push_mioi_biwt;
  input dma_read_ctrl_Push_mioi_bdwt;
  output dma_read_ctrl_Push_mioi_bcwt;
  reg dma_read_ctrl_Push_mioi_bcwt;
  input dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dma_read_ctrl_Push_mioi_wen_comp = (~ dma_read_ctrl_Push_mioi_oswt) | dma_read_ctrl_Push_mioi_biwt
      | dma_read_ctrl_Push_mioi_bcwt;
  assign dma_read_ctrl_Push_mioi_m_index_rsc_dat = {(dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input[31:7])
      , (~ dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_pff) , (~ dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_pff)
      , (~ dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_pff) , (~ dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_pff)
      , (~ dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_pff) , (~ dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_pff)
      , (~ dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_pff)};
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_read_ctrl_Push_mioi_bcwt <= ~((~(dma_read_ctrl_Push_mioi_bcwt | dma_read_ctrl_Push_mioi_biwt))
          | dma_read_ctrl_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl
    (
  load_input_wen, dma_read_ctrl_Push_mioi_oswt, dma_read_ctrl_Push_mioi_biwt, dma_read_ctrl_Push_mioi_bdwt,
      dma_read_ctrl_Push_mioi_bcwt, dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld,
      dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_pff, dma_read_ctrl_Push_mioi_oswt_pff
);
  input load_input_wen;
  input dma_read_ctrl_Push_mioi_oswt;
  output dma_read_ctrl_Push_mioi_biwt;
  output dma_read_ctrl_Push_mioi_bdwt;
  input dma_read_ctrl_Push_mioi_bcwt;
  input dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  output dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_pff;
  input dma_read_ctrl_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dma_read_ctrl_Push_mioi_bdwt = dma_read_ctrl_Push_mioi_oswt & load_input_wen;
  assign dma_read_ctrl_Push_mioi_biwt = dma_read_ctrl_Push_mioi_oswt & (~ dma_read_ctrl_Push_mioi_bcwt)
      & dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  assign dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_pff = dma_read_ctrl_Push_mioi_oswt_pff
      & load_input_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_config_accelerator_config_accelerator_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_config_accelerator_config_accelerator_fsm (
  clk, rst, fsm_output, CONFIG_LOOP_C_0_tr0
);
  input clk;
  input rst;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;
  input CONFIG_LOOP_C_0_tr0;


  // FSM State Type Declaration for esp_acc_softmax_softmax_config_accelerator_config_accelerator_fsm_1
  parameter
    config_accelerator_rlp_C_0 = 2'd0,
    CONFIG_LOOP_C_0 = 2'd1,
    CONFIG_DONE_LOOP_C_0 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_softmax_softmax_config_accelerator_config_accelerator_fsm_1
    case (state_var)
      CONFIG_LOOP_C_0 : begin
        fsm_output = 3'b010;
        if ( CONFIG_LOOP_C_0_tr0 ) begin
          state_var_NS = CONFIG_LOOP_C_0;
        end
        else begin
          state_var_NS = CONFIG_DONE_LOOP_C_0;
        end
      end
      CONFIG_DONE_LOOP_C_0 : begin
        fsm_output = 3'b100;
        state_var_NS = CONFIG_DONE_LOOP_C_0;
      end
      // config_accelerator_rlp_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = CONFIG_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= config_accelerator_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_req_obj
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_req_obj (
  clk, rst, plm_out_cns_req_vz, store_output_wen, plm_out_cns_req_obj_oswt, plm_out_cns_req_obj_wen_comp
);
  input clk;
  input rst;
  input plm_out_cns_req_vz;
  input store_output_wen;
  input plm_out_cns_req_obj_oswt;
  output plm_out_cns_req_obj_wen_comp;


  // Interconnect Declarations
  wire plm_out_cns_req_obj_vd;
  wire plm_out_cns_req_obj_biwt;
  wire plm_out_cns_req_obj_bdwt;
  wire plm_out_cns_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_mgc_in_sync_v2 #(.valid(32'sd1)) plm_out_cns_req_obj (
      .vd(plm_out_cns_req_obj_vd),
      .vz(plm_out_cns_req_vz)
    );
  esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl
      softmax_store_output_store_output_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl_inst
      (
      .store_output_wen(store_output_wen),
      .plm_out_cns_req_obj_oswt(plm_out_cns_req_obj_oswt),
      .plm_out_cns_req_obj_vd(plm_out_cns_req_obj_vd),
      .plm_out_cns_req_obj_biwt(plm_out_cns_req_obj_biwt),
      .plm_out_cns_req_obj_bdwt(plm_out_cns_req_obj_bdwt),
      .plm_out_cns_req_obj_bcwt(plm_out_cns_req_obj_bcwt)
    );
  esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_req_obj_plm_out_cns_req_wait_dp
      softmax_store_output_store_output_plm_out_cns_req_obj_plm_out_cns_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_req_obj_oswt(plm_out_cns_req_obj_oswt),
      .plm_out_cns_req_obj_wen_comp(plm_out_cns_req_obj_wen_comp),
      .plm_out_cns_req_obj_biwt(plm_out_cns_req_obj_biwt),
      .plm_out_cns_req_obj_bdwt(plm_out_cns_req_obj_bdwt),
      .plm_out_cns_req_obj_bcwt(plm_out_cns_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_rls_obj
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_rls_obj (
  plm_out_cns_rls_lz, store_output_wten, plm_out_cns_rls_obj_iswt0
);
  output plm_out_cns_rls_lz;
  input store_output_wten;
  input plm_out_cns_rls_obj_iswt0;


  // Interconnect Declarations
  wire plm_out_cns_rls_obj_ld_store_output_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_mgc_io_sync_v2 #(.valid(32'sd0)) plm_out_cns_rls_obj (
      .ld(plm_out_cns_rls_obj_ld_store_output_sct),
      .lz(plm_out_cns_rls_lz)
    );
  esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl
      softmax_store_output_store_output_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl_inst
      (
      .store_output_wten(store_output_wten),
      .plm_out_cns_rls_obj_iswt0(plm_out_cns_rls_obj_iswt0),
      .plm_out_cns_rls_obj_ld_store_output_sct(plm_out_cns_rls_obj_ld_store_output_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_1
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_1 (
  clk, rst, plm_out_cnsi_q_d, plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d, store_output_wen,
      store_output_wten, plm_out_cnsi_oswt, plm_out_cnsi_q_d_mxwt, plm_out_cnsi_oswt_pff
);
  input clk;
  input rst;
  input [31:0] plm_out_cnsi_q_d;
  output plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d;
  input store_output_wen;
  input store_output_wten;
  input plm_out_cnsi_oswt;
  output [31:0] plm_out_cnsi_q_d_mxwt;
  input plm_out_cnsi_oswt_pff;


  // Interconnect Declarations
  wire plm_out_cnsi_biwt;
  wire plm_out_cnsi_bdwt;
  wire plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_store_output_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_1_plm_out_cns_wait_ctrl
      softmax_store_output_store_output_plm_out_cnsi_1_plm_out_cns_wait_ctrl_inst
      (
      .store_output_wen(store_output_wen),
      .store_output_wten(store_output_wten),
      .plm_out_cnsi_oswt(plm_out_cnsi_oswt),
      .plm_out_cnsi_biwt(plm_out_cnsi_biwt),
      .plm_out_cnsi_bdwt(plm_out_cnsi_bdwt),
      .plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_store_output_sct(plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_store_output_sct),
      .plm_out_cnsi_oswt_pff(plm_out_cnsi_oswt_pff)
    );
  esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_1_plm_out_cns_wait_dp
      softmax_store_output_store_output_plm_out_cnsi_1_plm_out_cns_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_out_cnsi_q_d(plm_out_cnsi_q_d),
      .plm_out_cnsi_q_d_mxwt(plm_out_cnsi_q_d_mxwt),
      .plm_out_cnsi_biwt(plm_out_cnsi_biwt),
      .plm_out_cnsi_bdwt(plm_out_cnsi_bdwt)
    );
  assign plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d = plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_store_output_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi
    (
  clk, rst, dma_write_chnl_val, dma_write_chnl_rdy, dma_write_chnl_msg, store_output_wen,
      dma_write_chnl_Push_mioi_oswt, dma_write_chnl_Push_mioi_wen_comp, dma_write_chnl_Push_mioi_m_rsc_dat_store_output,
      dma_write_chnl_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;
  input store_output_wen;
  input dma_write_chnl_Push_mioi_oswt;
  output dma_write_chnl_Push_mioi_wen_comp;
  input [63:0] dma_write_chnl_Push_mioi_m_rsc_dat_store_output;
  input dma_write_chnl_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire [63:0] dma_write_chnl_Push_mioi_m_rsc_dat;
  wire dma_write_chnl_Push_mioi_biwt;
  wire dma_write_chnl_Push_mioi_bdwt;
  wire dma_write_chnl_Push_mioi_bcwt;
  wire dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld;
  wire dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [63:0] nl_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp_inst_dma_write_chnl_Push_mioi_m_rsc_dat_store_output;
  assign nl_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp_inst_dma_write_chnl_Push_mioi_m_rsc_dat_store_output
      = {32'b11011110101011011011111011101111 , (dma_write_chnl_Push_mioi_m_rsc_dat_store_output[31:0])};
  esp_acc_softmax_Connections_OutBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Push
      dma_write_chnl_Push_mioi (
      .this_val(dma_write_chnl_val),
      .this_rdy(dma_write_chnl_rdy),
      .this_msg(dma_write_chnl_msg),
      .m_rsc_dat(dma_write_chnl_Push_mioi_m_rsc_dat),
      .ccs_ccore_start_rsc_dat(dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_iff),
      .ccs_ccore_done_sync_vld(dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl
      softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl_inst
      (
      .store_output_wen(store_output_wen),
      .dma_write_chnl_Push_mioi_oswt(dma_write_chnl_Push_mioi_oswt),
      .dma_write_chnl_Push_mioi_biwt(dma_write_chnl_Push_mioi_biwt),
      .dma_write_chnl_Push_mioi_bdwt(dma_write_chnl_Push_mioi_bdwt),
      .dma_write_chnl_Push_mioi_bcwt(dma_write_chnl_Push_mioi_bcwt),
      .dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld(dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld),
      .dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff(dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_iff),
      .dma_write_chnl_Push_mioi_oswt_pff(dma_write_chnl_Push_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp
      softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_chnl_Push_mioi_oswt(dma_write_chnl_Push_mioi_oswt),
      .dma_write_chnl_Push_mioi_wen_comp(dma_write_chnl_Push_mioi_wen_comp),
      .dma_write_chnl_Push_mioi_m_rsc_dat_store_output(nl_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp_inst_dma_write_chnl_Push_mioi_m_rsc_dat_store_output[63:0]),
      .dma_write_chnl_Push_mioi_m_rsc_dat(dma_write_chnl_Push_mioi_m_rsc_dat),
      .dma_write_chnl_Push_mioi_biwt(dma_write_chnl_Push_mioi_biwt),
      .dma_write_chnl_Push_mioi_bdwt(dma_write_chnl_Push_mioi_bdwt),
      .dma_write_chnl_Push_mioi_bcwt(dma_write_chnl_Push_mioi_bcwt),
      .dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff(dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi
    (
  clk, rst, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg, store_output_wen,
      dma_write_ctrl_Push_mioi_oswt, dma_write_ctrl_Push_mioi_wen_comp, dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output,
      dma_write_ctrl_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  input store_output_wen;
  input dma_write_ctrl_Push_mioi_oswt;
  output dma_write_ctrl_Push_mioi_wen_comp;
  input [31:0] dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output;
  input dma_write_ctrl_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire [31:0] dma_write_ctrl_Push_mioi_m_index_rsc_dat;
  wire dma_write_ctrl_Push_mioi_biwt;
  wire dma_write_ctrl_Push_mioi_bdwt;
  wire dma_write_ctrl_Push_mioi_bcwt;
  wire dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  wire dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output;
  assign nl_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output
      = {(dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output[31:7]) , 7'b0000000};
  esp_acc_softmax_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push  dma_write_ctrl_Push_mioi
      (
      .this_val(dma_write_ctrl_val),
      .this_rdy(dma_write_ctrl_rdy),
      .this_msg(dma_write_ctrl_msg),
      .m_index_rsc_dat(dma_write_ctrl_Push_mioi_m_index_rsc_dat),
      .ccs_ccore_start_rsc_dat(dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_iff),
      .ccs_ccore_done_sync_vld(dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl
      softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl_inst
      (
      .store_output_wen(store_output_wen),
      .dma_write_ctrl_Push_mioi_oswt(dma_write_ctrl_Push_mioi_oswt),
      .dma_write_ctrl_Push_mioi_biwt(dma_write_ctrl_Push_mioi_biwt),
      .dma_write_ctrl_Push_mioi_bdwt(dma_write_ctrl_Push_mioi_bdwt),
      .dma_write_ctrl_Push_mioi_bcwt(dma_write_ctrl_Push_mioi_bcwt),
      .dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld(dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_pff(dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_iff),
      .dma_write_ctrl_Push_mioi_oswt_pff(dma_write_ctrl_Push_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp
      softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_ctrl_Push_mioi_oswt(dma_write_ctrl_Push_mioi_oswt),
      .dma_write_ctrl_Push_mioi_wen_comp(dma_write_ctrl_Push_mioi_wen_comp),
      .dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output(nl_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output[31:0]),
      .dma_write_ctrl_Push_mioi_m_index_rsc_dat(dma_write_ctrl_Push_mioi_m_index_rsc_dat),
      .dma_write_ctrl_Push_mioi_biwt(dma_write_ctrl_Push_mioi_biwt),
      .dma_write_ctrl_Push_mioi_bdwt(dma_write_ctrl_Push_mioi_bdwt),
      .dma_write_ctrl_Push_mioi_bcwt(dma_write_ctrl_Push_mioi_bcwt),
      .dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_pff(dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output_sct_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_output_ready_ack_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_output_ready_ack_mioi (
  clk, rst, output_ready_req_req, output_ready_ack_ack, store_output_wen, output_ready_ack_mioi_oswt,
      output_ready_ack_mioi_wen_comp, output_ready_ack_mioi_oswt_pff
);
  input clk;
  input rst;
  input output_ready_req_req;
  output output_ready_ack_ack;
  input store_output_wen;
  input output_ready_ack_mioi_oswt;
  output output_ready_ack_mioi_wen_comp;
  input output_ready_ack_mioi_oswt_pff;


  // Interconnect Declarations
  wire output_ready_ack_mioi_biwt;
  wire output_ready_ack_mioi_bdwt;
  wire output_ready_ack_mioi_bcwt;
  wire output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_output_sct;
  wire output_ready_ack_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_handshake_t_ack  output_ready_ack_mioi (
      .this_req_req(output_ready_req_req),
      .this_ack_ack(output_ready_ack_ack),
      .ccs_ccore_start_rsc_dat(output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_output_sct),
      .ccs_ccore_done_sync_vld(output_ready_ack_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_store_output_store_output_output_ready_ack_mioi_output_ready_ack_mio_wait_ctrl
      softmax_store_output_store_output_output_ready_ack_mioi_output_ready_ack_mio_wait_ctrl_inst
      (
      .store_output_wen(store_output_wen),
      .output_ready_ack_mioi_oswt(output_ready_ack_mioi_oswt),
      .output_ready_ack_mioi_biwt(output_ready_ack_mioi_biwt),
      .output_ready_ack_mioi_bdwt(output_ready_ack_mioi_bdwt),
      .output_ready_ack_mioi_bcwt(output_ready_ack_mioi_bcwt),
      .output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_output_sct(output_ready_ack_mioi_ccs_ccore_start_rsc_dat_store_output_sct),
      .output_ready_ack_mioi_ccs_ccore_done_sync_vld(output_ready_ack_mioi_ccs_ccore_done_sync_vld),
      .output_ready_ack_mioi_oswt_pff(output_ready_ack_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_store_output_store_output_output_ready_ack_mioi_output_ready_ack_mio_wait_dp
      softmax_store_output_store_output_output_ready_ack_mioi_output_ready_ack_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .output_ready_ack_mioi_oswt(output_ready_ack_mioi_oswt),
      .output_ready_ack_mioi_wen_comp(output_ready_ack_mioi_wen_comp),
      .output_ready_ack_mioi_biwt(output_ready_ack_mioi_biwt),
      .output_ready_ack_mioi_bdwt(output_ready_ack_mioi_bdwt),
      .output_ready_ack_mioi_bcwt(output_ready_ack_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_req_obj
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_req_obj
    (
  clk, rst, plm_out_cns_req_vz, compute_kernel_wen, plm_out_cns_req_obj_oswt, plm_out_cns_req_obj_wen_comp
);
  input clk;
  input rst;
  input plm_out_cns_req_vz;
  input compute_kernel_wen;
  input plm_out_cns_req_obj_oswt;
  output plm_out_cns_req_obj_wen_comp;


  // Interconnect Declarations
  wire plm_out_cns_req_obj_vd;
  wire plm_out_cns_req_obj_biwt;
  wire plm_out_cns_req_obj_bdwt;
  wire plm_out_cns_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_mgc_in_sync_v2 #(.valid(32'sd1)) plm_out_cns_req_obj (
      .vd(plm_out_cns_req_obj_vd),
      .vz(plm_out_cns_req_vz)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl
      softmax_compute_kernel_compute_kernel_plm_out_cns_req_obj_plm_out_cns_req_wait_ctrl_inst
      (
      .compute_kernel_wen(compute_kernel_wen),
      .plm_out_cns_req_obj_oswt(plm_out_cns_req_obj_oswt),
      .plm_out_cns_req_obj_vd(plm_out_cns_req_obj_vd),
      .plm_out_cns_req_obj_biwt(plm_out_cns_req_obj_biwt),
      .plm_out_cns_req_obj_bdwt(plm_out_cns_req_obj_bdwt),
      .plm_out_cns_req_obj_bcwt(plm_out_cns_req_obj_bcwt)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_req_obj_plm_out_cns_req_wait_dp
      softmax_compute_kernel_compute_kernel_plm_out_cns_req_obj_plm_out_cns_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_req_obj_oswt(plm_out_cns_req_obj_oswt),
      .plm_out_cns_req_obj_wen_comp(plm_out_cns_req_obj_wen_comp),
      .plm_out_cns_req_obj_biwt(plm_out_cns_req_obj_biwt),
      .plm_out_cns_req_obj_bdwt(plm_out_cns_req_obj_bdwt),
      .plm_out_cns_req_obj_bcwt(plm_out_cns_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_req_obj
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_req_obj (
  clk, rst, plm_in_cns_req_vz, compute_kernel_wen, plm_in_cns_req_obj_oswt, plm_in_cns_req_obj_wen_comp
);
  input clk;
  input rst;
  input plm_in_cns_req_vz;
  input compute_kernel_wen;
  input plm_in_cns_req_obj_oswt;
  output plm_in_cns_req_obj_wen_comp;


  // Interconnect Declarations
  wire plm_in_cns_req_obj_vd;
  wire plm_in_cns_req_obj_biwt;
  wire plm_in_cns_req_obj_bdwt;
  wire plm_in_cns_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_mgc_in_sync_v2 #(.valid(32'sd1)) plm_in_cns_req_obj (
      .vd(plm_in_cns_req_obj_vd),
      .vz(plm_in_cns_req_vz)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl
      softmax_compute_kernel_compute_kernel_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl_inst
      (
      .compute_kernel_wen(compute_kernel_wen),
      .plm_in_cns_req_obj_oswt(plm_in_cns_req_obj_oswt),
      .plm_in_cns_req_obj_vd(plm_in_cns_req_obj_vd),
      .plm_in_cns_req_obj_biwt(plm_in_cns_req_obj_biwt),
      .plm_in_cns_req_obj_bdwt(plm_in_cns_req_obj_bdwt),
      .plm_in_cns_req_obj_bcwt(plm_in_cns_req_obj_bcwt)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_req_obj_plm_in_cns_req_wait_dp
      softmax_compute_kernel_compute_kernel_plm_in_cns_req_obj_plm_in_cns_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_req_obj_oswt(plm_in_cns_req_obj_oswt),
      .plm_in_cns_req_obj_wen_comp(plm_in_cns_req_obj_wen_comp),
      .plm_in_cns_req_obj_biwt(plm_in_cns_req_obj_biwt),
      .plm_in_cns_req_obj_bdwt(plm_in_cns_req_obj_bdwt),
      .plm_in_cns_req_obj_bcwt(plm_in_cns_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_rls_obj
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_rls_obj (
  plm_in_cns_rls_lz, compute_kernel_wten, plm_in_cns_rls_obj_iswt0
);
  output plm_in_cns_rls_lz;
  input compute_kernel_wten;
  input plm_in_cns_rls_obj_iswt0;


  // Interconnect Declarations
  wire plm_in_cns_rls_obj_ld_compute_kernel_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_mgc_io_sync_v2 #(.valid(32'sd0)) plm_in_cns_rls_obj (
      .ld(plm_in_cns_rls_obj_ld_compute_kernel_sct),
      .lz(plm_in_cns_rls_lz)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl
      softmax_compute_kernel_compute_kernel_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl_inst
      (
      .compute_kernel_wten(compute_kernel_wten),
      .plm_in_cns_rls_obj_iswt0(plm_in_cns_rls_obj_iswt0),
      .plm_in_cns_rls_obj_ld_compute_kernel_sct(plm_in_cns_rls_obj_ld_compute_kernel_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_rls_obj
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_rls_obj
    (
  plm_out_cns_rls_lz, compute_kernel_wten, plm_out_cns_rls_obj_iswt0
);
  output plm_out_cns_rls_lz;
  input compute_kernel_wten;
  input plm_out_cns_rls_obj_iswt0;


  // Interconnect Declarations
  wire plm_out_cns_rls_obj_ld_compute_kernel_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_mgc_io_sync_v2 #(.valid(32'sd0)) plm_out_cns_rls_obj (
      .ld(plm_out_cns_rls_obj_ld_compute_kernel_sct),
      .lz(plm_out_cns_rls_lz)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl
      softmax_compute_kernel_compute_kernel_plm_out_cns_rls_obj_plm_out_cns_rls_wait_ctrl_inst
      (
      .compute_kernel_wten(compute_kernel_wten),
      .plm_out_cns_rls_obj_iswt0(plm_out_cns_rls_obj_iswt0),
      .plm_out_cns_rls_obj_ld_compute_kernel_sct(plm_out_cns_rls_obj_ld_compute_kernel_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi_1
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi_1 (
  plm_out_cnsi_we_d_pff, plm_out_cnsi_iswt0_pff, compute_kernel_wten_pff
);
  output plm_out_cnsi_we_d_pff;
  input plm_out_cnsi_iswt0_pff;
  input compute_kernel_wten_pff;


  // Interconnect Declarations
  wire plm_out_cnsi_we_d_compute_kernel_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi_1_plm_out_cns_wait_ctrl
      softmax_compute_kernel_compute_kernel_plm_out_cnsi_1_plm_out_cns_wait_ctrl_inst
      (
      .plm_out_cnsi_we_d_compute_kernel_sct_pff(plm_out_cnsi_we_d_compute_kernel_sct_iff),
      .plm_out_cnsi_iswt0_pff(plm_out_cnsi_iswt0_pff),
      .compute_kernel_wten_pff(compute_kernel_wten_pff)
    );
  assign plm_out_cnsi_we_d_pff = plm_out_cnsi_we_d_compute_kernel_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_1
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_1 (
  clk, rst, plm_in_cnsi_q_d, plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d, compute_kernel_wen,
      compute_kernel_wten, plm_in_cnsi_oswt, plm_in_cnsi_q_d_mxwt, plm_in_cnsi_oswt_pff
);
  input clk;
  input rst;
  input [31:0] plm_in_cnsi_q_d;
  output plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d;
  input compute_kernel_wen;
  input compute_kernel_wten;
  input plm_in_cnsi_oswt;
  output [31:0] plm_in_cnsi_q_d_mxwt;
  input plm_in_cnsi_oswt_pff;


  // Interconnect Declarations
  wire plm_in_cnsi_biwt;
  wire plm_in_cnsi_bdwt;
  wire plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_compute_kernel_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_1_plm_in_cns_wait_ctrl
      softmax_compute_kernel_compute_kernel_plm_in_cnsi_1_plm_in_cns_wait_ctrl_inst
      (
      .compute_kernel_wen(compute_kernel_wen),
      .compute_kernel_wten(compute_kernel_wten),
      .plm_in_cnsi_oswt(plm_in_cnsi_oswt),
      .plm_in_cnsi_biwt(plm_in_cnsi_biwt),
      .plm_in_cnsi_bdwt(plm_in_cnsi_bdwt),
      .plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_compute_kernel_sct(plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_compute_kernel_sct),
      .plm_in_cnsi_oswt_pff(plm_in_cnsi_oswt_pff)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_1_plm_in_cns_wait_dp
      softmax_compute_kernel_compute_kernel_plm_in_cnsi_1_plm_in_cns_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cnsi_q_d(plm_in_cnsi_q_d),
      .plm_in_cnsi_q_d_mxwt(plm_in_cnsi_q_d_mxwt),
      .plm_in_cnsi_biwt(plm_in_cnsi_biwt),
      .plm_in_cnsi_bdwt(plm_in_cnsi_bdwt)
    );
  assign plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d = plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_compute_kernel_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_req_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_req_mioi
    (
  clk, rst, output_ready_req_req, output_ready_ack_ack, compute_kernel_wen, output_ready_req_mioi_oswt,
      output_ready_req_mioi_wen_comp, output_ready_req_mioi_oswt_pff
);
  input clk;
  input rst;
  output output_ready_req_req;
  input output_ready_ack_ack;
  input compute_kernel_wen;
  input output_ready_req_mioi_oswt;
  output output_ready_req_mioi_wen_comp;
  input output_ready_req_mioi_oswt_pff;


  // Interconnect Declarations
  wire output_ready_req_mioi_biwt;
  wire output_ready_req_mioi_bdwt;
  wire output_ready_req_mioi_bcwt;
  wire output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct;
  wire output_ready_req_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_handshake_t_req  output_ready_req_mioi (
      .this_req_req(output_ready_req_req),
      .this_ack_ack(output_ready_ack_ack),
      .ccs_ccore_start_rsc_dat(output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct),
      .ccs_ccore_done_sync_vld(output_ready_req_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_req_mioi_output_ready_req_mio_wait_ctrl
      softmax_compute_kernel_compute_kernel_output_ready_req_mioi_output_ready_req_mio_wait_ctrl_inst
      (
      .compute_kernel_wen(compute_kernel_wen),
      .output_ready_req_mioi_oswt(output_ready_req_mioi_oswt),
      .output_ready_req_mioi_biwt(output_ready_req_mioi_biwt),
      .output_ready_req_mioi_bdwt(output_ready_req_mioi_bdwt),
      .output_ready_req_mioi_bcwt(output_ready_req_mioi_bcwt),
      .output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct(output_ready_req_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct),
      .output_ready_req_mioi_ccs_ccore_done_sync_vld(output_ready_req_mioi_ccs_ccore_done_sync_vld),
      .output_ready_req_mioi_oswt_pff(output_ready_req_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_req_mioi_output_ready_req_mio_wait_dp
      softmax_compute_kernel_compute_kernel_output_ready_req_mioi_output_ready_req_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .output_ready_req_mioi_oswt(output_ready_req_mioi_oswt),
      .output_ready_req_mioi_wen_comp(output_ready_req_mioi_wen_comp),
      .output_ready_req_mioi_biwt(output_ready_req_mioi_biwt),
      .output_ready_req_mioi_bdwt(output_ready_req_mioi_bdwt),
      .output_ready_req_mioi_bcwt(output_ready_req_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_ack_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_ack_mioi
    (
  clk, rst, input_ready_req_req, input_ready_ack_ack, compute_kernel_wen, input_ready_ack_mioi_oswt,
      input_ready_ack_mioi_wen_comp, input_ready_ack_mioi_oswt_pff
);
  input clk;
  input rst;
  input input_ready_req_req;
  output input_ready_ack_ack;
  input compute_kernel_wen;
  input input_ready_ack_mioi_oswt;
  output input_ready_ack_mioi_wen_comp;
  input input_ready_ack_mioi_oswt_pff;


  // Interconnect Declarations
  wire input_ready_ack_mioi_biwt;
  wire input_ready_ack_mioi_bdwt;
  wire input_ready_ack_mioi_bcwt;
  wire input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct;
  wire input_ready_ack_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_handshake_t_ack  input_ready_ack_mioi (
      .this_req_req(input_ready_req_req),
      .this_ack_ack(input_ready_ack_ack),
      .ccs_ccore_start_rsc_dat(input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct),
      .ccs_ccore_done_sync_vld(input_ready_ack_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_ack_mioi_input_ready_ack_mio_wait_ctrl
      softmax_compute_kernel_compute_kernel_input_ready_ack_mioi_input_ready_ack_mio_wait_ctrl_inst
      (
      .compute_kernel_wen(compute_kernel_wen),
      .input_ready_ack_mioi_oswt(input_ready_ack_mioi_oswt),
      .input_ready_ack_mioi_biwt(input_ready_ack_mioi_biwt),
      .input_ready_ack_mioi_bdwt(input_ready_ack_mioi_bdwt),
      .input_ready_ack_mioi_bcwt(input_ready_ack_mioi_bcwt),
      .input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct(input_ready_ack_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct),
      .input_ready_ack_mioi_ccs_ccore_done_sync_vld(input_ready_ack_mioi_ccs_ccore_done_sync_vld),
      .input_ready_ack_mioi_oswt_pff(input_ready_ack_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_ack_mioi_input_ready_ack_mio_wait_dp
      softmax_compute_kernel_compute_kernel_input_ready_ack_mioi_input_ready_ack_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_ready_ack_mioi_oswt(input_ready_ack_mioi_oswt),
      .input_ready_ack_mioi_wen_comp(input_ready_ack_mioi_wen_comp),
      .input_ready_ack_mioi_biwt(input_ready_ack_mioi_biwt),
      .input_ready_ack_mioi_bdwt(input_ready_ack_mioi_bdwt),
      .input_ready_ack_mioi_bcwt(input_ready_ack_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_req_obj
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_req_obj (
  clk, rst, plm_in_cns_req_vz, load_input_wen, plm_in_cns_req_obj_oswt, plm_in_cns_req_obj_wen_comp
);
  input clk;
  input rst;
  input plm_in_cns_req_vz;
  input load_input_wen;
  input plm_in_cns_req_obj_oswt;
  output plm_in_cns_req_obj_wen_comp;


  // Interconnect Declarations
  wire plm_in_cns_req_obj_vd;
  wire plm_in_cns_req_obj_biwt;
  wire plm_in_cns_req_obj_bdwt;
  wire plm_in_cns_req_obj_bcwt;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_mgc_in_sync_v2 #(.valid(32'sd1)) plm_in_cns_req_obj (
      .vd(plm_in_cns_req_obj_vd),
      .vz(plm_in_cns_req_vz)
    );
  esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl
      softmax_load_input_load_input_plm_in_cns_req_obj_plm_in_cns_req_wait_ctrl_inst
      (
      .load_input_wen(load_input_wen),
      .plm_in_cns_req_obj_oswt(plm_in_cns_req_obj_oswt),
      .plm_in_cns_req_obj_vd(plm_in_cns_req_obj_vd),
      .plm_in_cns_req_obj_biwt(plm_in_cns_req_obj_biwt),
      .plm_in_cns_req_obj_bdwt(plm_in_cns_req_obj_bdwt),
      .plm_in_cns_req_obj_bcwt(plm_in_cns_req_obj_bcwt)
    );
  esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_req_obj_plm_in_cns_req_wait_dp
      softmax_load_input_load_input_plm_in_cns_req_obj_plm_in_cns_req_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_req_obj_oswt(plm_in_cns_req_obj_oswt),
      .plm_in_cns_req_obj_wen_comp(plm_in_cns_req_obj_wen_comp),
      .plm_in_cns_req_obj_biwt(plm_in_cns_req_obj_biwt),
      .plm_in_cns_req_obj_bdwt(plm_in_cns_req_obj_bdwt),
      .plm_in_cns_req_obj_bcwt(plm_in_cns_req_obj_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_rls_obj
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_rls_obj (
  plm_in_cns_rls_lz, load_input_wten, plm_in_cns_rls_obj_iswt0
);
  output plm_in_cns_rls_lz;
  input load_input_wten;
  input plm_in_cns_rls_obj_iswt0;


  // Interconnect Declarations
  wire plm_in_cns_rls_obj_ld_load_input_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_mgc_io_sync_v2 #(.valid(32'sd0)) plm_in_cns_rls_obj (
      .ld(plm_in_cns_rls_obj_ld_load_input_sct),
      .lz(plm_in_cns_rls_lz)
    );
  esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl
      softmax_load_input_load_input_plm_in_cns_rls_obj_plm_in_cns_rls_wait_ctrl_inst
      (
      .load_input_wten(load_input_wten),
      .plm_in_cns_rls_obj_iswt0(plm_in_cns_rls_obj_iswt0),
      .plm_in_cns_rls_obj_ld_load_input_sct(plm_in_cns_rls_obj_ld_load_input_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi_1
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi_1 (
  plm_in_cnsi_we_d_pff, plm_in_cnsi_iswt0_pff, load_input_wten_pff
);
  output plm_in_cnsi_we_d_pff;
  input plm_in_cnsi_iswt0_pff;
  input load_input_wten_pff;


  // Interconnect Declarations
  wire plm_in_cnsi_we_d_load_input_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi_1_plm_in_cns_wait_ctrl
      softmax_load_input_load_input_plm_in_cnsi_1_plm_in_cns_wait_ctrl_inst (
      .plm_in_cnsi_we_d_load_input_sct_pff(plm_in_cnsi_we_d_load_input_sct_iff),
      .plm_in_cnsi_iswt0_pff(plm_in_cnsi_iswt0_pff),
      .load_input_wten_pff(load_input_wten_pff)
    );
  assign plm_in_cnsi_we_d_pff = plm_in_cnsi_we_d_load_input_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_input_ready_req_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_input_ready_req_mioi (
  clk, rst, input_ready_req_req, input_ready_ack_ack, load_input_wen, input_ready_req_mioi_oswt,
      input_ready_req_mioi_wen_comp, input_ready_req_mioi_oswt_pff
);
  input clk;
  input rst;
  output input_ready_req_req;
  input input_ready_ack_ack;
  input load_input_wen;
  input input_ready_req_mioi_oswt;
  output input_ready_req_mioi_wen_comp;
  input input_ready_req_mioi_oswt_pff;


  // Interconnect Declarations
  wire input_ready_req_mioi_biwt;
  wire input_ready_req_mioi_bdwt;
  wire input_ready_req_mioi_bcwt;
  wire input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_input_sct;
  wire input_ready_req_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_handshake_t_req  input_ready_req_mioi (
      .this_req_req(input_ready_req_req),
      .this_ack_ack(input_ready_ack_ack),
      .ccs_ccore_start_rsc_dat(input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_input_sct),
      .ccs_ccore_done_sync_vld(input_ready_req_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_load_input_load_input_input_ready_req_mioi_input_ready_req_mio_wait_ctrl
      softmax_load_input_load_input_input_ready_req_mioi_input_ready_req_mio_wait_ctrl_inst
      (
      .load_input_wen(load_input_wen),
      .input_ready_req_mioi_oswt(input_ready_req_mioi_oswt),
      .input_ready_req_mioi_biwt(input_ready_req_mioi_biwt),
      .input_ready_req_mioi_bdwt(input_ready_req_mioi_bdwt),
      .input_ready_req_mioi_bcwt(input_ready_req_mioi_bcwt),
      .input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_input_sct(input_ready_req_mioi_ccs_ccore_start_rsc_dat_load_input_sct),
      .input_ready_req_mioi_ccs_ccore_done_sync_vld(input_ready_req_mioi_ccs_ccore_done_sync_vld),
      .input_ready_req_mioi_oswt_pff(input_ready_req_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_load_input_load_input_input_ready_req_mioi_input_ready_req_mio_wait_dp
      softmax_load_input_load_input_input_ready_req_mioi_input_ready_req_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_ready_req_mioi_oswt(input_ready_req_mioi_oswt),
      .input_ready_req_mioi_wen_comp(input_ready_req_mioi_wen_comp),
      .input_ready_req_mioi_biwt(input_ready_req_mioi_biwt),
      .input_ready_req_mioi_bdwt(input_ready_req_mioi_bdwt),
      .input_ready_req_mioi_bcwt(input_ready_req_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi (
  clk, rst, dma_read_chnl_val, dma_read_chnl_rdy, dma_read_chnl_msg, load_input_wen,
      dma_read_chnl_Pop_mioi_oswt, dma_read_chnl_Pop_mioi_wen_comp, dma_read_chnl_Pop_mioi_return_rsc_z_mxwt,
      dma_read_chnl_Pop_mioi_oswt_pff
);
  input clk;
  input rst;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  input load_input_wen;
  input dma_read_chnl_Pop_mioi_oswt;
  output dma_read_chnl_Pop_mioi_wen_comp;
  output [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt;
  input dma_read_chnl_Pop_mioi_oswt_pff;


  // Interconnect Declarations
  wire [63:0] dma_read_chnl_Pop_mioi_return_rsc_z;
  wire dma_read_chnl_Pop_mioi_biwt;
  wire dma_read_chnl_Pop_mioi_bdwt;
  wire dma_read_chnl_Pop_mioi_bcwt;
  wire dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct;
  wire dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld;
  wire [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_Connections_InBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Pop
      dma_read_chnl_Pop_mioi (
      .this_val(dma_read_chnl_val),
      .this_rdy(dma_read_chnl_rdy),
      .this_msg(dma_read_chnl_msg),
      .return_rsc_z(dma_read_chnl_Pop_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct),
      .ccs_ccore_done_sync_vld(dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl
      softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl_inst
      (
      .load_input_wen(load_input_wen),
      .dma_read_chnl_Pop_mioi_oswt(dma_read_chnl_Pop_mioi_oswt),
      .dma_read_chnl_Pop_mioi_biwt(dma_read_chnl_Pop_mioi_biwt),
      .dma_read_chnl_Pop_mioi_bdwt(dma_read_chnl_Pop_mioi_bdwt),
      .dma_read_chnl_Pop_mioi_bcwt(dma_read_chnl_Pop_mioi_bcwt),
      .dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct(dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct),
      .dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld(dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld),
      .dma_read_chnl_Pop_mioi_oswt_pff(dma_read_chnl_Pop_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp
      softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_chnl_Pop_mioi_oswt(dma_read_chnl_Pop_mioi_oswt),
      .dma_read_chnl_Pop_mioi_wen_comp(dma_read_chnl_Pop_mioi_wen_comp),
      .dma_read_chnl_Pop_mioi_return_rsc_z_mxwt(dma_read_chnl_Pop_mioi_return_rsc_z_mxwt_pconst),
      .dma_read_chnl_Pop_mioi_return_rsc_z(dma_read_chnl_Pop_mioi_return_rsc_z),
      .dma_read_chnl_Pop_mioi_biwt(dma_read_chnl_Pop_mioi_biwt),
      .dma_read_chnl_Pop_mioi_bdwt(dma_read_chnl_Pop_mioi_bdwt),
      .dma_read_chnl_Pop_mioi_bcwt(dma_read_chnl_Pop_mioi_bcwt)
    );
  assign dma_read_chnl_Pop_mioi_return_rsc_z_mxwt = dma_read_chnl_Pop_mioi_return_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi (
  clk, rst, dma_read_ctrl_val, dma_read_ctrl_rdy, dma_read_ctrl_msg, load_input_wen,
      dma_read_ctrl_Push_mioi_oswt, dma_read_ctrl_Push_mioi_wen_comp, dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input,
      dma_read_ctrl_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  input load_input_wen;
  input dma_read_ctrl_Push_mioi_oswt;
  output dma_read_ctrl_Push_mioi_wen_comp;
  input [31:0] dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input;
  input dma_read_ctrl_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire [31:0] dma_read_ctrl_Push_mioi_m_index_rsc_dat;
  wire dma_read_ctrl_Push_mioi_biwt;
  wire dma_read_ctrl_Push_mioi_bdwt;
  wire dma_read_ctrl_Push_mioi_bcwt;
  wire dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  wire dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input;
  assign nl_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input
      = {(dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input[31:7]) , 7'b0000000};
  esp_acc_softmax_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push  dma_read_ctrl_Push_mioi
      (
      .this_val(dma_read_ctrl_val),
      .this_rdy(dma_read_ctrl_rdy),
      .this_msg(dma_read_ctrl_msg),
      .m_index_rsc_dat(dma_read_ctrl_Push_mioi_m_index_rsc_dat),
      .ccs_ccore_start_rsc_dat(dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_iff),
      .ccs_ccore_done_sync_vld(dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl
      softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl_inst
      (
      .load_input_wen(load_input_wen),
      .dma_read_ctrl_Push_mioi_oswt(dma_read_ctrl_Push_mioi_oswt),
      .dma_read_ctrl_Push_mioi_biwt(dma_read_ctrl_Push_mioi_biwt),
      .dma_read_ctrl_Push_mioi_bdwt(dma_read_ctrl_Push_mioi_bdwt),
      .dma_read_ctrl_Push_mioi_bcwt(dma_read_ctrl_Push_mioi_bcwt),
      .dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld(dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_pff(dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_iff),
      .dma_read_ctrl_Push_mioi_oswt_pff(dma_read_ctrl_Push_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp
      softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_ctrl_Push_mioi_oswt(dma_read_ctrl_Push_mioi_oswt),
      .dma_read_ctrl_Push_mioi_wen_comp(dma_read_ctrl_Push_mioi_wen_comp),
      .dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input(nl_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input[31:0]),
      .dma_read_ctrl_Push_mioi_m_index_rsc_dat(dma_read_ctrl_Push_mioi_m_index_rsc_dat),
      .dma_read_ctrl_Push_mioi_biwt(dma_read_ctrl_Push_mioi_biwt),
      .dma_read_ctrl_Push_mioi_bdwt(dma_read_ctrl_Push_mioi_bdwt),
      .dma_read_ctrl_Push_mioi_bcwt(dma_read_ctrl_Push_mioi_bcwt),
      .dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_pff(dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input_sct_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_config_accelerator
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_config_accelerator (
  clk, rst, conf_done, done
);
  input clk;
  input rst;
  input conf_done;
  output done;
  reg done;


  // Interconnect Declarations
  wire [2:0] fsm_output;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_softmax_config_accelerator_config_accelerator_fsm_inst_CONFIG_LOOP_C_0_tr0;
  assign nl_softmax_config_accelerator_config_accelerator_fsm_inst_CONFIG_LOOP_C_0_tr0
      = ~ conf_done;
  esp_acc_softmax_softmax_config_accelerator_config_accelerator_fsm softmax_config_accelerator_config_accelerator_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .CONFIG_LOOP_C_0_tr0(nl_softmax_config_accelerator_config_accelerator_fsm_inst_CONFIG_LOOP_C_0_tr0[0:0])
    );
  always @(posedge clk) begin
    if ( ~ rst ) begin
      done <= 1'b0;
    end
    else if ( conf_done & (fsm_output[1]) ) begin
      done <= 1'b1;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output (
  clk, rst, conf_info, acc_done, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg,
      dma_write_chnl_val, dma_write_chnl_rdy, dma_write_chnl_msg, done, output_ready_req_req,
      output_ready_ack_ack, plm_out_cns_req_vz, plm_out_cns_rls_lz, plm_out_cnsi_q_d,
      plm_out_cnsi_radr_d, plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d
);
  input clk;
  input rst;
  input [31:0] conf_info;
  output acc_done;
  reg acc_done;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;
  input done;
  input output_ready_req_req;
  output output_ready_ack_ack;
  input plm_out_cns_req_vz;
  output plm_out_cns_rls_lz;
  input [31:0] plm_out_cnsi_q_d;
  output [6:0] plm_out_cnsi_radr_d;
  output plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations
  wire store_output_wen;
  wire store_output_wten;
  wire output_ready_ack_mioi_wen_comp;
  wire dma_write_ctrl_Push_mioi_wen_comp;
  wire dma_write_chnl_Push_mioi_wen_comp;
  wire [31:0] plm_out_cnsi_q_d_mxwt;
  wire plm_out_cns_req_obj_wen_comp;
  wire [6:0] fsm_output;
  wire [7:0] STORE_DATA_INNER_LOOP_acc_1_tmp;
  wire [8:0] nl_STORE_DATA_INNER_LOOP_acc_1_tmp;
  wire and_dcpl_12;
  reg exitL_exit_STORE_DATA_INNER_LOOP_sva;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_st_1;
  reg STORE_BATCH_LOOP_stage_0_1;
  reg exit_STORE_BATCH_LOOP_sva_1_st_1;
  reg STORE_BATCH_LOOP_stage_0_2;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3;
  reg STORE_BATCH_LOOP_stage_0_4;
  reg exit_STORE_BATCH_LOOP_lpi_1_dfm_st_2;
  reg reg_output_ready_ack_mioi_oswt_cse;
  reg reg_dma_write_ctrl_Push_mioi_oswt_cse;
  reg reg_dma_write_chnl_Push_mioi_oswt_cse;
  reg reg_plm_out_cnsi_oswt_cse;
  reg reg_plm_out_cns_rls_obj_iswt0_cse;
  reg reg_STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_7_1_itm_2_cse;
  wire plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_reg;
  wire and_31_rmff;
  wire and_21_rmff;
  wire and_23_rmff;
  wire and_27_rmff;
  reg [6:0] STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_6_0_itm_2;
  reg [24:0] STORE_BATCH_LOOP_asn_2_itm_1;
  reg [31:0] config_batch_sva;
  reg [24:0] offset_31_7_sva;
  reg [31:0] STORE_BATCH_LOOP_b_sva;
  reg STORE_BATCH_LOOP_stage_0_3;
  reg [6:0] STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_6_0_itm_1;
  wire [6:0] STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_6_0_itm_1_mx0;
  reg [6:0] STORE_DATA_INNER_LOOP_i_7_0_sva_1_6_0;
  wire offset_and_1_rgt;
  wire STORE_BATCH_LOOP_acc_itm_32_1;

  wire[31:0] STORE_BATCH_LOOP_b_mux_nl;
  wire[31:0] STORE_BATCH_LOOP_acc_2_nl;
  wire[32:0] nl_STORE_BATCH_LOOP_acc_2_nl;
  wire[0:0] STORE_BATCH_LOOP_b_and_nl;
  wire[24:0] STORE_BATCH_LOOP_acc_1_nl;
  wire[25:0] nl_STORE_BATCH_LOOP_acc_1_nl;
  wire[32:0] STORE_BATCH_LOOP_acc_nl;
  wire[33:0] nl_STORE_BATCH_LOOP_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output;
  assign nl_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output
      = {STORE_BATCH_LOOP_asn_2_itm_1 , 7'b0000000};
  wire [63:0] nl_softmax_store_output_store_output_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_m_rsc_dat_store_output;
  assign nl_softmax_store_output_store_output_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_m_rsc_dat_store_output
      = {32'b11011110101011011011111011101111 , plm_out_cnsi_q_d_mxwt};
  wire [0:0] nl_softmax_store_output_store_output_store_output_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  assign nl_softmax_store_output_store_output_store_output_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0
      = ~ done;
  wire [0:0] nl_softmax_store_output_store_output_store_output_fsm_inst_STORE_BATCH_LOOP_C_0_tr0;
  assign nl_softmax_store_output_store_output_store_output_fsm_inst_STORE_BATCH_LOOP_C_0_tr0
      = STORE_BATCH_LOOP_stage_0_3 | STORE_BATCH_LOOP_stage_0_4 | STORE_BATCH_LOOP_stage_0_2
      | STORE_BATCH_LOOP_stage_0_1;
  esp_acc_softmax_softmax_store_output_store_output_output_ready_ack_mioi softmax_store_output_store_output_output_ready_ack_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .output_ready_req_req(output_ready_req_req),
      .output_ready_ack_ack(output_ready_ack_ack),
      .store_output_wen(store_output_wen),
      .output_ready_ack_mioi_oswt(reg_output_ready_ack_mioi_oswt_cse),
      .output_ready_ack_mioi_wen_comp(output_ready_ack_mioi_wen_comp),
      .output_ready_ack_mioi_oswt_pff(and_21_rmff)
    );
  esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi softmax_store_output_store_output_dma_write_ctrl_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_ctrl_val(dma_write_ctrl_val),
      .dma_write_ctrl_rdy(dma_write_ctrl_rdy),
      .dma_write_ctrl_msg(dma_write_ctrl_msg),
      .store_output_wen(store_output_wen),
      .dma_write_ctrl_Push_mioi_oswt(reg_dma_write_ctrl_Push_mioi_oswt_cse),
      .dma_write_ctrl_Push_mioi_wen_comp(dma_write_ctrl_Push_mioi_wen_comp),
      .dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output(nl_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output[31:0]),
      .dma_write_ctrl_Push_mioi_oswt_pff(and_23_rmff)
    );
  esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi softmax_store_output_store_output_dma_write_chnl_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_chnl_val(dma_write_chnl_val),
      .dma_write_chnl_rdy(dma_write_chnl_rdy),
      .dma_write_chnl_msg(dma_write_chnl_msg),
      .store_output_wen(store_output_wen),
      .dma_write_chnl_Push_mioi_oswt(reg_dma_write_chnl_Push_mioi_oswt_cse),
      .dma_write_chnl_Push_mioi_wen_comp(dma_write_chnl_Push_mioi_wen_comp),
      .dma_write_chnl_Push_mioi_m_rsc_dat_store_output(nl_softmax_store_output_store_output_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_m_rsc_dat_store_output[63:0]),
      .dma_write_chnl_Push_mioi_oswt_pff(and_27_rmff)
    );
  esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_1 softmax_store_output_store_output_plm_out_cnsi_1_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cnsi_q_d(plm_out_cnsi_q_d),
      .plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d(plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_reg),
      .store_output_wen(store_output_wen),
      .store_output_wten(store_output_wten),
      .plm_out_cnsi_oswt(reg_plm_out_cnsi_oswt_cse),
      .plm_out_cnsi_q_d_mxwt(plm_out_cnsi_q_d_mxwt),
      .plm_out_cnsi_oswt_pff(and_31_rmff)
    );
  esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_rls_obj softmax_store_output_store_output_plm_out_cns_rls_obj_inst
      (
      .plm_out_cns_rls_lz(plm_out_cns_rls_lz),
      .store_output_wten(store_output_wten),
      .plm_out_cns_rls_obj_iswt0(reg_plm_out_cns_rls_obj_iswt0_cse)
    );
  esp_acc_softmax_softmax_store_output_store_output_plm_out_cns_req_obj softmax_store_output_store_output_plm_out_cns_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_req_vz(plm_out_cns_req_vz),
      .store_output_wen(store_output_wen),
      .plm_out_cns_req_obj_oswt(reg_dma_write_ctrl_Push_mioi_oswt_cse),
      .plm_out_cns_req_obj_wen_comp(plm_out_cns_req_obj_wen_comp)
    );
  esp_acc_softmax_softmax_store_output_store_output_staller softmax_store_output_store_output_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .store_output_wen(store_output_wen),
      .store_output_wten(store_output_wten),
      .output_ready_ack_mioi_wen_comp(output_ready_ack_mioi_wen_comp),
      .dma_write_ctrl_Push_mioi_wen_comp(dma_write_ctrl_Push_mioi_wen_comp),
      .dma_write_chnl_Push_mioi_wen_comp(dma_write_chnl_Push_mioi_wen_comp),
      .plm_out_cns_req_obj_wen_comp(plm_out_cns_req_obj_wen_comp)
    );
  esp_acc_softmax_softmax_store_output_store_output_store_output_fsm softmax_store_output_store_output_store_output_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .store_output_wen(store_output_wen),
      .fsm_output(fsm_output),
      .WAIT_FOR_CONFIG_LOOP_C_0_tr0(nl_softmax_store_output_store_output_store_output_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0[0:0]),
      .STORE_BATCH_LOOP_C_0_tr0(nl_softmax_store_output_store_output_store_output_fsm_inst_STORE_BATCH_LOOP_C_0_tr0[0:0])
    );
  assign and_21_rmff = exitL_exit_STORE_DATA_INNER_LOOP_sva & STORE_BATCH_LOOP_stage_0_1
      & STORE_BATCH_LOOP_acc_itm_32_1 & (fsm_output[1]);
  assign and_23_rmff = STORE_BATCH_LOOP_stage_0_2 & (~ exit_STORE_BATCH_LOOP_sva_1_st_1)
      & reg_STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_7_1_itm_2_cse
      & (fsm_output[1]);
  assign and_27_rmff = STORE_BATCH_LOOP_stage_0_4 & (~ exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3)
      & (fsm_output[1]);
  assign and_31_rmff = and_dcpl_12 & (fsm_output[1]);
  assign offset_and_1_rgt = exitL_exit_STORE_DATA_INNER_LOOP_sva & (fsm_output[1]);
  assign nl_STORE_BATCH_LOOP_acc_nl = ({1'b1 , STORE_BATCH_LOOP_b_sva}) + conv_u2u_32_33(~
      config_batch_sva) + 33'b000000000000000000000000000000001;
  assign STORE_BATCH_LOOP_acc_nl = nl_STORE_BATCH_LOOP_acc_nl[32:0];
  assign STORE_BATCH_LOOP_acc_itm_32_1 = readslicef_33_1_32(STORE_BATCH_LOOP_acc_nl);
  assign nl_STORE_DATA_INNER_LOOP_acc_1_tmp = conv_u2u_7_8(STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_6_0_itm_1_mx0)
      + 8'b00000001;
  assign STORE_DATA_INNER_LOOP_acc_1_tmp = nl_STORE_DATA_INNER_LOOP_acc_1_tmp[7:0];
  assign STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_6_0_itm_1_mx0 =
      MUX_v_7_2_2(STORE_DATA_INNER_LOOP_i_7_0_sva_1_6_0, (signext_7_1(~ STORE_BATCH_LOOP_acc_itm_32_1)),
      exitL_exit_STORE_DATA_INNER_LOOP_sva);
  assign and_dcpl_12 = STORE_BATCH_LOOP_stage_0_3 & (~ exit_STORE_BATCH_LOOP_lpi_1_dfm_st_2);
  assign plm_out_cnsi_radr_d = STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_6_0_itm_2;
  assign plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d = plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      acc_done <= 1'b0;
    end
    else if ( store_output_wen & ((fsm_output[5]) | (fsm_output[2])) ) begin
      acc_done <= ~ (fsm_output[5]);
    end
  end
  always @(posedge clk) begin
    if ( store_output_wen ) begin
      STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_6_0_itm_2 <= STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_6_0_itm_1;
      STORE_BATCH_LOOP_asn_2_itm_1 <= offset_31_7_sva;
      STORE_BATCH_LOOP_b_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          STORE_BATCH_LOOP_b_mux_nl, (fsm_output[1]));
      config_batch_sva <= MUX_v_32_2_2(conf_info, config_batch_sva, fsm_output[1]);
      STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_6_0_itm_1 <= STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_6_0_itm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_output_ready_ack_mioi_oswt_cse <= 1'b0;
      reg_dma_write_ctrl_Push_mioi_oswt_cse <= 1'b0;
      reg_dma_write_chnl_Push_mioi_oswt_cse <= 1'b0;
      reg_plm_out_cnsi_oswt_cse <= 1'b0;
      reg_plm_out_cns_rls_obj_iswt0_cse <= 1'b0;
      STORE_BATCH_LOOP_stage_0_1 <= 1'b0;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3 <= 1'b0;
      reg_STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_7_1_itm_2_cse <=
          1'b0;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_st_2 <= 1'b0;
      exit_STORE_BATCH_LOOP_sva_1_st_1 <= 1'b0;
      STORE_DATA_INNER_LOOP_i_7_0_sva_1_6_0 <= 7'b0000000;
      exitL_exit_STORE_DATA_INNER_LOOP_sva <= 1'b0;
      STORE_BATCH_LOOP_stage_0_2 <= 1'b0;
      STORE_BATCH_LOOP_stage_0_3 <= 1'b0;
      STORE_BATCH_LOOP_stage_0_4 <= 1'b0;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_st_1 <= 1'b0;
    end
    else if ( store_output_wen ) begin
      reg_output_ready_ack_mioi_oswt_cse <= and_21_rmff;
      reg_dma_write_ctrl_Push_mioi_oswt_cse <= and_23_rmff;
      reg_dma_write_chnl_Push_mioi_oswt_cse <= and_27_rmff;
      reg_plm_out_cnsi_oswt_cse <= and_31_rmff;
      reg_plm_out_cns_rls_obj_iswt0_cse <= and_dcpl_12 & reg_STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_7_1_itm_2_cse
          & (fsm_output[1]);
      STORE_BATCH_LOOP_stage_0_1 <= ~((~(STORE_BATCH_LOOP_stage_0_1 & ((~ exitL_exit_STORE_DATA_INNER_LOOP_sva)
          | STORE_BATCH_LOOP_acc_itm_32_1))) & (fsm_output[1]));
      exit_STORE_BATCH_LOOP_lpi_1_dfm_st_3 <= exit_STORE_BATCH_LOOP_lpi_1_dfm_st_2;
      reg_STORE_DATA_INNER_LOOP_i_slc_STORE_DATA_INNER_LOOP_i_7_0_7_1_itm_2_cse <=
          exitL_exit_STORE_DATA_INNER_LOOP_sva;
      exit_STORE_BATCH_LOOP_lpi_1_dfm_st_2 <= exit_STORE_BATCH_LOOP_lpi_1_dfm_st_1;
      exit_STORE_BATCH_LOOP_sva_1_st_1 <= ~ STORE_BATCH_LOOP_acc_itm_32_1;
      STORE_DATA_INNER_LOOP_i_7_0_sva_1_6_0 <= STORE_DATA_INNER_LOOP_acc_1_tmp[6:0];
      exitL_exit_STORE_DATA_INNER_LOOP_sva <= (STORE_DATA_INNER_LOOP_acc_1_tmp[7])
          | (~ (fsm_output[1]));
      STORE_BATCH_LOOP_stage_0_2 <= STORE_BATCH_LOOP_stage_0_1 & (fsm_output[1]);
      STORE_BATCH_LOOP_stage_0_3 <= STORE_BATCH_LOOP_stage_0_2 & (fsm_output[1]);
      STORE_BATCH_LOOP_stage_0_4 <= STORE_BATCH_LOOP_stage_0_3 & (fsm_output[1]);
      exit_STORE_BATCH_LOOP_lpi_1_dfm_st_1 <= (~ STORE_BATCH_LOOP_acc_itm_32_1) &
          exitL_exit_STORE_DATA_INNER_LOOP_sva;
    end
  end
  always @(posedge clk) begin
    if ( store_output_wen & ((~ (fsm_output[1])) | offset_and_1_rgt) ) begin
      offset_31_7_sva <= MUX_v_25_2_2((conf_info[24:0]), STORE_BATCH_LOOP_acc_1_nl,
          offset_and_1_rgt);
    end
  end
  assign nl_STORE_BATCH_LOOP_acc_2_nl = STORE_BATCH_LOOP_b_sva + 32'b00000000000000000000000000000001;
  assign STORE_BATCH_LOOP_acc_2_nl = nl_STORE_BATCH_LOOP_acc_2_nl[31:0];
  assign STORE_BATCH_LOOP_b_and_nl = (STORE_DATA_INNER_LOOP_acc_1_tmp[7]) & (fsm_output[1]);
  assign STORE_BATCH_LOOP_b_mux_nl = MUX_v_32_2_2(STORE_BATCH_LOOP_b_sva, STORE_BATCH_LOOP_acc_2_nl,
      STORE_BATCH_LOOP_b_and_nl);
  assign nl_STORE_BATCH_LOOP_acc_1_nl = offset_31_7_sva + 25'b0000000000000000000000001;
  assign STORE_BATCH_LOOP_acc_1_nl = nl_STORE_BATCH_LOOP_acc_1_nl[24:0];

  function automatic [24:0] MUX_v_25_2_2;
    input [24:0] input_0;
    input [24:0] input_1;
    input [0:0] sel;
    reg [24:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_25_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input [0:0] vector;
  begin
    signext_7_1= {{6{vector[0]}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [32:0] conv_u2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_33 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel (
  clk, rst, conf_info, done, input_ready_req_req, input_ready_ack_ack, output_ready_req_req,
      output_ready_ack_ack, plm_in_cns_req_vz, plm_in_cns_rls_lz, plm_out_cns_req_vz,
      plm_out_cns_rls_lz, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      plm_in_cnsi_q_d, plm_in_cnsi_radr_d, plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d,
      plm_out_cnsi_d_d, plm_out_cnsi_wadr_d, CALC_SOFTMAX_LOOP_mul_cmp_b, CALC_SOFTMAX_LOOP_mul_cmp_z,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d_pff,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff,
      plm_out_cnsi_we_d_pff
);
  input clk;
  input rst;
  input [31:0] conf_info;
  input done;
  input input_ready_req_req;
  output input_ready_ack_ack;
  output output_ready_req_req;
  input output_ready_ack_ack;
  input plm_in_cns_req_vz;
  output plm_in_cns_rls_lz;
  input plm_out_cns_req_vz;
  output plm_out_cns_rls_lz;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d;
  output [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  input [31:0] plm_in_cnsi_q_d;
  output [6:0] plm_in_cnsi_radr_d;
  output plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d;
  output [31:0] plm_out_cnsi_d_d;
  output [6:0] plm_out_cnsi_wadr_d;
  output [93:0] CALC_SOFTMAX_LOOP_mul_cmp_b;
  input [94:0] CALC_SOFTMAX_LOOP_mul_cmp_z;
  output [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d_pff;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff;
  output plm_out_cnsi_we_d_pff;


  // Interconnect Declarations
  wire compute_kernel_wen;
  wire compute_kernel_wten;
  wire input_ready_ack_mioi_wen_comp;
  wire output_ready_req_mioi_wen_comp;
  wire [31:0] plm_in_cnsi_q_d_mxwt;
  wire plm_in_cns_req_obj_wen_comp;
  wire plm_out_cns_req_obj_wen_comp;
  wire [2:0] fsm_output;
  wire [7:0] CALC_SOFTMAX_LOOP_acc_1_tmp;
  wire [8:0] nl_CALC_SOFTMAX_LOOP_acc_1_tmp;
  wire [73:0] SUM_EXP_LOOP_acc_1_tmp;
  wire [74:0] nl_SUM_EXP_LOOP_acc_1_tmp;
  wire [7:0] SUM_EXP_LOOP_acc_2_tmp;
  wire [8:0] nl_SUM_EXP_LOOP_acc_2_tmp;
  wire [7:0] CALC_EXP_LOOP_acc_1_tmp;
  wire [8:0] nl_CALC_EXP_LOOP_acc_1_tmp;
  wire and_dcpl_50;
  wire and_dcpl_60;
  wire and_dcpl_63;
  wire or_dcpl_12;
  wire and_dcpl_77;
  reg exitL_exit_CALC_SOFTMAX_LOOP_sva;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1_1;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1;
  wire CALC_SOFTMAX_LOOP_and_4_ssc_1;
  wire CALC_SOFTMAX_LOOP_and_5_ssc_1;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0_mx0;
  wire CALC_SOFTMAX_LOOP_equal_tmp_2;
  wire CALC_SOFTMAX_LOOP_or_tmp_1;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1_mx0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_7;
  reg CALC_SOFTMAX_LOOP_asn_itm_6;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1;
  reg COMPUTE_BATCH_LOOP_asn_2_itm_4;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_3;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_2;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0;
  reg CALC_SOFTMAX_LOOP_and_10_itm_4;
  reg CALC_SOFTMAX_LOOP_asn_itm_2;
  reg COMPUTE_BATCH_LOOP_stage_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_6;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1;
  reg CALC_SOFTMAX_LOOP_asn_itm_5;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1;
  reg COMPUTE_BATCH_LOOP_asn_2_itm_5;
  reg CALC_SOFTMAX_LOOP_asn_itm_4;
  reg CALC_SOFTMAX_LOOP_asn_itm_1;
  reg CALC_SOFTMAX_LOOP_asn_itm_3;
  reg COMPUTE_BATCH_LOOP_stage_0_10;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9;
  reg exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_8;
  reg CALC_EXP_LOOP_and_svs_st_2;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_st_1;
  reg COMPUTE_BATCH_LOOP_stage_0_2;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_st_7;
  reg COMPUTE_BATCH_LOOP_stage_0_8;
  reg CALC_SOFTMAX_LOOP_asn_itm_7;
  reg CALC_SOFTMAX_LOOP_and_10_itm_5;
  reg COMPUTE_BATCH_LOOP_stage_0_6;
  reg CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_4;
  reg COMPUTE_BATCH_LOOP_stage_0_5;
  reg CALC_EXP_LOOP_and_svs_st_4;
  wire or_14_tmp;
  reg reg_input_ready_ack_mioi_oswt_cse;
  reg reg_output_ready_req_mioi_oswt_cse;
  reg reg_plm_in_cnsi_oswt_cse;
  reg reg_plm_out_cns_rls_obj_iswt0_cse;
  reg reg_plm_in_cns_rls_obj_iswt0_cse;
  reg reg_plm_in_cns_req_obj_oswt_cse;
  reg reg_plm_out_cns_req_obj_oswt_cse;
  wire ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_and_cse;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_and_cse;
  wire and_76_cse;
  wire plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_reg;
  wire and_167_rmff;
  wire plm_out_cnsi_we_d_iff;
  wire and_163_rmff;
  wire and_165_rmff;
  reg [6:0] CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_2_6_0;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_8;
  reg [93:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1;
  reg [66:0] operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1;
  reg [6:0] CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_2;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_3;
  wire [73:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_mx1;
  wire [93:0] operator_94_21_false_AC_TRN_AC_WRAP_rshift_itm;
  wire [66:0] operator_67_47_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [72:0] operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm;
  reg [73:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1;
  reg [31:0] config_batch_sva;
  reg [31:0] COMPUTE_BATCH_LOOP_b_sva;
  reg COMPUTE_BATCH_LOOP_stage_0_3;
  reg COMPUTE_BATCH_LOOP_stage_0_4;
  reg COMPUTE_BATCH_LOOP_stage_0_7;
  reg COMPUTE_BATCH_LOOP_stage_0_9;
  reg [10:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm;
  wire [11:0] nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm;
  reg [9:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_9_0_itm;
  reg [7:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm;
  wire [8:0] nl_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_2;
  reg [73:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_1_1;
  reg [6:0] CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_1;
  reg ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_itm_1;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_5;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_6;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_7;
  reg CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_1;
  reg CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_2;
  reg CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_3;
  reg CALC_SOFTMAX_LOOP_and_10_itm_1;
  reg CALC_SOFTMAX_LOOP_and_10_itm_2;
  reg CALC_SOFTMAX_LOOP_and_10_itm_3;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_st_4;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_st_5;
  reg exit_COMPUTE_BATCH_LOOP_sva_1_st_6;
  reg CALC_EXP_LOOP_and_svs_st_1;
  reg CALC_EXP_LOOP_and_svs_st_3;
  reg CALC_EXP_LOOP_and_svs_st_5;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_6;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_7;
  reg [6:0] CALC_EXP_LOOP_i_7_0_lpi_1_6_0;
  reg [6:0] SUM_EXP_LOOP_i_7_0_lpi_1_6_0;
  reg [6:0] CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_1_6_0;
  wire [6:0] CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_1_6_0_mx0;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire [18:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire signed [19:0] nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire [6:0] libraries_leading_sign_74_0_cfd8a2a1b60025d53198d215150438e7bf24_1;
  wire COMPUTE_BATCH_LOOP_acc_itm_32_1;
  wire [18:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1;

  wire[93:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_or_nl;
  wire[0:0] or_8_nl;
  wire[0:0] or_nl;
  wire[31:0] COMPUTE_BATCH_LOOP_b_mux_nl;
  wire[31:0] COMPUTE_BATCH_LOOP_acc_1_nl;
  wire[32:0] nl_COMPUTE_BATCH_LOOP_acc_1_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_b_and_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_and_14_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_and_15_nl;
  wire[9:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl;
  wire[32:0] COMPUTE_BATCH_LOOP_acc_nl;
  wire[33:0] nl_COMPUTE_BATCH_LOOP_acc_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_24_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_2_nl;
  wire[0:0] and_74_nl;
  wire[0:0] and_75_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_and_5_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_and_6_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_nl;
  wire[2:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_1_nl;
  wire[46:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl;
  wire signed [47:0] nl_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl;
  wire[6:0] CALC_SOFTMAX_LOOP_mux_29_nl;
  wire[7:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [73:0] nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_a;
  assign nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_a = {ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm
      , ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_9_0_itm
      , 53'b00000000000000000000000000000000000000000000000000000};
  wire[10:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[2:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_2_nl;
  wire[6:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_3_nl;
  wire [20:0] nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_2_nl
      = MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1[11:10]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_3_nl
      = MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1[11:10]);
  assign nl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:10])
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_2_nl
      , 1'b1 , ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_3_nl});
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a = {ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , (ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[9:0])};
  wire [6:0] nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_s = ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1[18:12];
  wire [72:0] nl_operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg_a = SUM_EXP_LOOP_acc_1_tmp[72:0];
  wire [0:0] nl_softmax_compute_kernel_compute_kernel_plm_out_cnsi_1_inst_plm_out_cnsi_iswt0_pff;
  assign nl_softmax_compute_kernel_compute_kernel_plm_out_cnsi_1_inst_plm_out_cnsi_iswt0_pff
      = and_dcpl_63 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0) & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1
      & (fsm_output[1]);
  wire [0:0] nl_softmax_compute_kernel_compute_kernel_plm_out_cnsi_1_inst_compute_kernel_wten_pff;
  assign nl_softmax_compute_kernel_compute_kernel_plm_out_cnsi_1_inst_compute_kernel_wten_pff
      = ~ compute_kernel_wen;
  wire [0:0] nl_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  assign nl_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0
      = ~ done;
  wire [0:0] nl_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_inst_COMPUTE_BATCH_LOOP_C_0_tr0;
  assign nl_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_inst_COMPUTE_BATCH_LOOP_C_0_tr0
      = COMPUTE_BATCH_LOOP_stage_0 | COMPUTE_BATCH_LOOP_stage_0_2 | COMPUTE_BATCH_LOOP_stage_0_3
      | COMPUTE_BATCH_LOOP_stage_0_4 | COMPUTE_BATCH_LOOP_stage_0_5 | COMPUTE_BATCH_LOOP_stage_0_6
      | COMPUTE_BATCH_LOOP_stage_0_7 | COMPUTE_BATCH_LOOP_stage_0_8 | COMPUTE_BATCH_LOOP_stage_0_9
      | COMPUTE_BATCH_LOOP_stage_0_10;
  esp_acc_softmax_mgc_shift_br_v5 #(.width_a(32'sd74),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd94)) operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_a[73:0]),
      .s(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm),
      .z(operator_94_21_false_AC_TRN_AC_WRAP_rshift_itm)
    );
  esp_acc_softmax_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd67)) operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_s[6:0]),
      .z(operator_67_47_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  esp_acc_softmax_mgc_shift_l_v5 #(.width_a(32'sd73),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd73)) operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg_a[72:0]),
      .s(libraries_leading_sign_74_0_cfd8a2a1b60025d53198d215150438e7bf24_1),
      .z(operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  esp_acc_softmax_leading_sign_74_0  leading_sign_74_0_rg (
      .mantissa(SUM_EXP_LOOP_acc_1_tmp),
      .rtn(libraries_leading_sign_74_0_cfd8a2a1b60025d53198d215150438e7bf24_1)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_ack_mioi softmax_compute_kernel_compute_kernel_input_ready_ack_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .input_ready_req_req(input_ready_req_req),
      .input_ready_ack_ack(input_ready_ack_ack),
      .compute_kernel_wen(compute_kernel_wen),
      .input_ready_ack_mioi_oswt(reg_input_ready_ack_mioi_oswt_cse),
      .input_ready_ack_mioi_wen_comp(input_ready_ack_mioi_wen_comp),
      .input_ready_ack_mioi_oswt_pff(and_163_rmff)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_req_mioi softmax_compute_kernel_compute_kernel_output_ready_req_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .output_ready_req_req(output_ready_req_req),
      .output_ready_ack_ack(output_ready_ack_ack),
      .compute_kernel_wen(compute_kernel_wen),
      .output_ready_req_mioi_oswt(reg_output_ready_req_mioi_oswt_cse),
      .output_ready_req_mioi_wen_comp(output_ready_req_mioi_wen_comp),
      .output_ready_req_mioi_oswt_pff(and_165_rmff)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_1 softmax_compute_kernel_compute_kernel_plm_in_cnsi_1_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cnsi_q_d(plm_in_cnsi_q_d),
      .plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d(plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_reg),
      .compute_kernel_wen(compute_kernel_wen),
      .compute_kernel_wten(compute_kernel_wten),
      .plm_in_cnsi_oswt(reg_plm_in_cnsi_oswt_cse),
      .plm_in_cnsi_q_d_mxwt(plm_in_cnsi_q_d_mxwt),
      .plm_in_cnsi_oswt_pff(and_167_rmff)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi_1 softmax_compute_kernel_compute_kernel_plm_out_cnsi_1_inst
      (
      .plm_out_cnsi_we_d_pff(plm_out_cnsi_we_d_iff),
      .plm_out_cnsi_iswt0_pff(nl_softmax_compute_kernel_compute_kernel_plm_out_cnsi_1_inst_plm_out_cnsi_iswt0_pff[0:0]),
      .compute_kernel_wten_pff(nl_softmax_compute_kernel_compute_kernel_plm_out_cnsi_1_inst_compute_kernel_wten_pff[0:0])
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_rls_obj softmax_compute_kernel_compute_kernel_plm_out_cns_rls_obj_inst
      (
      .plm_out_cns_rls_lz(plm_out_cns_rls_lz),
      .compute_kernel_wten(compute_kernel_wten),
      .plm_out_cns_rls_obj_iswt0(reg_plm_out_cns_rls_obj_iswt0_cse)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_rls_obj softmax_compute_kernel_compute_kernel_plm_in_cns_rls_obj_inst
      (
      .plm_in_cns_rls_lz(plm_in_cns_rls_lz),
      .compute_kernel_wten(compute_kernel_wten),
      .plm_in_cns_rls_obj_iswt0(reg_plm_in_cns_rls_obj_iswt0_cse)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cns_req_obj softmax_compute_kernel_compute_kernel_plm_in_cns_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_req_vz(plm_in_cns_req_vz),
      .compute_kernel_wen(compute_kernel_wen),
      .plm_in_cns_req_obj_oswt(reg_plm_in_cns_req_obj_oswt_cse),
      .plm_in_cns_req_obj_wen_comp(plm_in_cns_req_obj_wen_comp)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cns_req_obj softmax_compute_kernel_compute_kernel_plm_out_cns_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_req_vz(plm_out_cns_req_vz),
      .compute_kernel_wen(compute_kernel_wen),
      .plm_out_cns_req_obj_oswt(reg_plm_out_cns_req_obj_oswt_cse),
      .plm_out_cns_req_obj_wen_comp(plm_out_cns_req_obj_wen_comp)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_staller softmax_compute_kernel_compute_kernel_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .compute_kernel_wen(compute_kernel_wen),
      .compute_kernel_wten(compute_kernel_wten),
      .input_ready_ack_mioi_wen_comp(input_ready_ack_mioi_wen_comp),
      .output_ready_req_mioi_wen_comp(output_ready_req_mioi_wen_comp),
      .plm_in_cns_req_obj_wen_comp(plm_in_cns_req_obj_wen_comp),
      .plm_out_cns_req_obj_wen_comp(plm_out_cns_req_obj_wen_comp)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_compute_kernel_fsm softmax_compute_kernel_compute_kernel_compute_kernel_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .compute_kernel_wen(compute_kernel_wen),
      .fsm_output(fsm_output),
      .WAIT_FOR_CONFIG_LOOP_C_0_tr0(nl_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0[0:0]),
      .COMPUTE_BATCH_LOOP_C_0_tr0(nl_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_inst_COMPUTE_BATCH_LOOP_C_0_tr0[0:0])
    );
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d
      = compute_kernel_wen;
  assign and_163_rmff = COMPUTE_BATCH_LOOP_acc_itm_32_1 & exitL_exit_CALC_SOFTMAX_LOOP_sva
      & COMPUTE_BATCH_LOOP_stage_0 & (fsm_output[1]);
  assign and_165_rmff = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0)
      & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9) & COMPUTE_BATCH_LOOP_stage_0_10
      & CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9 & (fsm_output[1]);
  assign and_167_rmff = and_dcpl_60 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1)
      & (fsm_output[1]);
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_and_cse
      = compute_kernel_wen & (fsm_output[1]);
  assign and_76_cse = (CALC_EXP_LOOP_acc_1_tmp[7]) & (SUM_EXP_LOOP_acc_2_tmp[7]);
  assign or_14_tmp = and_dcpl_77 | and_76_cse;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_and_cse = compute_kernel_wen
      & (~(((SUM_EXP_LOOP_acc_1_tmp==74'b00000000000000000000000000000000000000000000000000000000000000000000000000))
      | or_dcpl_12 | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1 | (~ CALC_EXP_LOOP_and_svs_st_4)
      | (~ (fsm_output[1]))));
  assign nl_SUM_EXP_LOOP_acc_1_tmp = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_1_1
      + conv_u2u_67_74(operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1);
  assign SUM_EXP_LOOP_acc_1_tmp = nl_SUM_EXP_LOOP_acc_1_tmp[73:0];
  assign nl_COMPUTE_BATCH_LOOP_acc_nl = ({1'b1 , COMPUTE_BATCH_LOOP_b_sva}) + conv_u2u_32_33(~
      config_batch_sva) + 33'b000000000000000000000000000000001;
  assign COMPUTE_BATCH_LOOP_acc_nl = nl_COMPUTE_BATCH_LOOP_acc_nl[32:0];
  assign COMPUTE_BATCH_LOOP_acc_itm_32_1 = readslicef_33_1_32(COMPUTE_BATCH_LOOP_acc_nl);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_2_nl = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1_mx0
      & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0_mx0;
  assign CALC_SOFTMAX_LOOP_mux_24_nl = MUX_s_1_2_2((~ (CALC_SOFTMAX_LOOP_acc_1_tmp[7])),
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1, CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_2_nl);
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1_1 = (CALC_SOFTMAX_LOOP_mux_24_nl
      & (~ CALC_SOFTMAX_LOOP_and_4_ssc_1)) | CALC_SOFTMAX_LOOP_and_5_ssc_1;
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0_1 = (lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0_mx0
      & (~(CALC_SOFTMAX_LOOP_and_5_ssc_1 | CALC_SOFTMAX_LOOP_equal_tmp_2))) | CALC_SOFTMAX_LOOP_and_4_ssc_1;
  assign and_74_nl = and_dcpl_50 & CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_4;
  assign and_75_nl = and_dcpl_50 & (~ CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_4);
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_mx1
      = MUX1HOT_v_74_3_2(SUM_EXP_LOOP_acc_1_tmp, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_1_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1,
      {and_74_nl , and_75_nl , or_dcpl_12});
  assign COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_and_5_nl = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1
      & (~ COMPUTE_BATCH_LOOP_acc_itm_32_1);
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1_mx0 = MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1,
      COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_and_5_nl, exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_and_6_nl = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0
      & (~ COMPUTE_BATCH_LOOP_acc_itm_32_1);
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0_mx0 = MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0,
      COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_and_6_nl, exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_1_6_0_mx0 = MUX_v_7_2_2(CALC_EXP_LOOP_i_7_0_lpi_1_6_0,
      (signext_7_1(~ COMPUTE_BATCH_LOOP_acc_itm_32_1)), exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign CALC_SOFTMAX_LOOP_or_tmp_1 = (lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0_mx0
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1_mx0)) | (~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1_mx0
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0_mx0));
  assign CALC_SOFTMAX_LOOP_and_5_ssc_1 = and_76_cse & CALC_SOFTMAX_LOOP_or_tmp_1;
  assign nl_CALC_SOFTMAX_LOOP_acc_1_tmp = conv_u2u_7_8(CALC_EXP_LOOP_i_7_0_lpi_1_6_0)
      + 8'b00000001;
  assign CALC_SOFTMAX_LOOP_acc_1_tmp = nl_CALC_SOFTMAX_LOOP_acc_1_tmp[7:0];
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1[11:10]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_1_nl
      = MUX_v_3_4_2(3'b010, 3'b110, 3'b001, 3'b101, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1[11:10]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = conv_u2u_19_19(({ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_nl
      , 1'b0 , ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_1_nl})
      * (ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1[9:0]));
  assign nl_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl
      = $signed((plm_in_cnsi_q_d_mxwt)) * $signed(16'b0101110001010101);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl
      = nl_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl[46:0];
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1
      = readslicef_47_19_28(ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl);
  assign CALC_SOFTMAX_LOOP_equal_tmp_2 = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1_mx0
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0_mx0);
  assign nl_CALC_EXP_LOOP_acc_1_tmp = conv_u2u_7_8(CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_1_6_0_mx0)
      + 8'b00000001;
  assign CALC_EXP_LOOP_acc_1_tmp = nl_CALC_EXP_LOOP_acc_1_tmp[7:0];
  assign CALC_SOFTMAX_LOOP_mux_29_nl = MUX_v_7_2_2(SUM_EXP_LOOP_i_7_0_lpi_1_6_0,
      (signext_7_1(~ COMPUTE_BATCH_LOOP_acc_itm_32_1)), exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign nl_SUM_EXP_LOOP_acc_2_tmp = conv_u2u_7_8(CALC_SOFTMAX_LOOP_mux_29_nl) +
      8'b00000001;
  assign SUM_EXP_LOOP_acc_2_tmp = nl_SUM_EXP_LOOP_acc_2_tmp[7:0];
  assign CALC_SOFTMAX_LOOP_and_4_ssc_1 = (~ and_76_cse) & CALC_SOFTMAX_LOOP_or_tmp_1;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_3_nl
      = MUX_v_8_8_2(8'b00011100, 8'b01001011, 8'b01101100, 8'b10000100, 8'b10010111,
      8'b10100110, 8'b10110011, 8'b10111100, operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm[72:70]);
  assign nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = $signed(({1'b1 , ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_3_nl}))
      * $signed(conv_u2s_10_11(operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm[69:60]));
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:0];
  assign and_dcpl_50 = COMPUTE_BATCH_LOOP_stage_0_5 & (~ COMPUTE_BATCH_LOOP_asn_2_itm_4);
  assign and_dcpl_60 = COMPUTE_BATCH_LOOP_stage_0_3 & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_2);
  assign and_dcpl_63 = COMPUTE_BATCH_LOOP_stage_0_9 & (~ exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8);
  assign or_dcpl_12 = (~ COMPUTE_BATCH_LOOP_stage_0_5) | COMPUTE_BATCH_LOOP_asn_2_itm_4;
  assign and_dcpl_77 = (~ exitL_exit_CALC_SOFTMAX_LOOP_sva) & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1;
  assign CALC_SOFTMAX_LOOP_mul_cmp_b = ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d
      = operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d_pff
      = CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_2;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff
      = and_dcpl_50 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1) & (fsm_output[1]);
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = and_dcpl_50 & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0)
      & (fsm_output[1]);
  assign plm_in_cnsi_radr_d = CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_2_6_0;
  assign plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d = plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d_reg;
  assign plm_out_cnsi_d_d = CALC_SOFTMAX_LOOP_mul_cmp_z[94:63];
  assign plm_out_cnsi_wadr_d = CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_8;
  assign plm_out_cnsi_we_d_pff = plm_out_cnsi_we_d_iff;
  always @(posedge clk) begin
    if ( compute_kernel_wen ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_8 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_7;
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_1_1
          <= MUX_v_74_2_2(({{73{exit_COMPUTE_BATCH_LOOP_sva_1_3}}, exit_COMPUTE_BATCH_LOOP_sva_1_3}),
          ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_mx1,
          or_nl);
      operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1 <= operator_67_47_false_AC_TRN_AC_WRAP_lshift_itm;
      CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_2 <= CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_1;
      CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_2_6_0 <= CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_1_6_0;
      COMPUTE_BATCH_LOOP_b_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          COMPUTE_BATCH_LOOP_b_mux_nl, (fsm_output[1]));
      config_batch_sva <= MUX_v_32_2_2(conf_info, config_batch_sva, fsm_output[1]);
      SUM_EXP_LOOP_i_7_0_lpi_1_6_0 <= SUM_EXP_LOOP_acc_2_tmp[6:0];
      CALC_EXP_LOOP_i_7_0_lpi_1_6_0 <= MUX1HOT_v_7_3_2((CALC_EXP_LOOP_acc_1_tmp[6:0]),
          (signext_7_1(~ and_76_cse)), (CALC_SOFTMAX_LOOP_acc_1_tmp[6:0]), {(~ or_14_tmp)
          , CALC_SOFTMAX_LOOP_and_14_nl , CALC_SOFTMAX_LOOP_and_15_nl});
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_7 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_6;
      CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_1 <= CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_2_6_0;
      CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_1_6_0 <= CALC_EXP_LOOP_i_7_0_lpi_1_dfm_1_1_6_0_mx0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_6 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_5;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_1_itm_5 <= CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_input_ready_ack_mioi_oswt_cse <= 1'b0;
      reg_output_ready_req_mioi_oswt_cse <= 1'b0;
      reg_plm_in_cnsi_oswt_cse <= 1'b0;
      reg_plm_out_cns_rls_obj_iswt0_cse <= 1'b0;
      reg_plm_in_cns_rls_obj_iswt0_cse <= 1'b0;
      reg_plm_in_cns_req_obj_oswt_cse <= 1'b0;
      reg_plm_out_cns_req_obj_oswt_cse <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_8 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_7 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_7 <= 1'b0;
      CALC_EXP_LOOP_and_svs_st_5 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_0 <= 1'b0;
      COMPUTE_BATCH_LOOP_asn_2_itm_5 <= 1'b0;
      CALC_EXP_LOOP_and_svs_st_4 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0 <= 1'b0;
      COMPUTE_BATCH_LOOP_asn_2_itm_4 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_3 <= 1'b0;
      CALC_EXP_LOOP_and_svs_st_2 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_2 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_1 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0 <= 1'b0;
      exitL_exit_CALC_SOFTMAX_LOOP_sva <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_2 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_3 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_4 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_5 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_6 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_7 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_8 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_9 <= 1'b0;
      COMPUTE_BATCH_LOOP_stage_0_10 <= 1'b0;
      ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_itm_1
          <= 1'b0;
      CALC_SOFTMAX_LOOP_and_10_itm_5 <= 1'b0;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_4 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_sva_1_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_7 <= 1'b0;
      CALC_EXP_LOOP_and_svs_st_1 <= 1'b0;
      CALC_EXP_LOOP_and_svs_st_3 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_1 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_7 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_6 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_6 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_6 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_6 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_5 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_5 <= 1'b0;
      CALC_SOFTMAX_LOOP_and_10_itm_4 <= 1'b0;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_3 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_sva_1_2 <= 1'b0;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_4 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_4 <= 1'b0;
      CALC_SOFTMAX_LOOP_and_10_itm_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_and_10_itm_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_and_10_itm_1 <= 1'b0;
    end
    else if ( compute_kernel_wen ) begin
      reg_input_ready_ack_mioi_oswt_cse <= and_163_rmff;
      reg_output_ready_req_mioi_oswt_cse <= and_165_rmff;
      reg_plm_in_cnsi_oswt_cse <= and_167_rmff;
      reg_plm_out_cns_rls_obj_iswt0_cse <= and_dcpl_63 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0)
          & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1 & CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_8
          & (fsm_output[1]);
      reg_plm_in_cns_rls_obj_iswt0_cse <= and_dcpl_60 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1)
          & CALC_EXP_LOOP_and_svs_st_2 & (fsm_output[1]);
      reg_plm_in_cns_req_obj_oswt_cse <= COMPUTE_BATCH_LOOP_stage_0_2 & CALC_SOFTMAX_LOOP_asn_itm_1
          & (~ exit_COMPUTE_BATCH_LOOP_sva_1_st_1) & (fsm_output[1]);
      reg_plm_out_cns_req_obj_oswt_cse <= COMPUTE_BATCH_LOOP_stage_0_8 & CALC_SOFTMAX_LOOP_asn_itm_7
          & (~ exit_COMPUTE_BATCH_LOOP_sva_1_st_7) & (fsm_output[1]);
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_9 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_8;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_9_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_9 <= exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_8 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_7;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_8_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_8 <= exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_7;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_7 <= exit_COMPUTE_BATCH_LOOP_sva_1_st_6;
      CALC_SOFTMAX_LOOP_asn_itm_7 <= CALC_SOFTMAX_LOOP_asn_itm_6;
      CALC_EXP_LOOP_and_svs_st_5 <= CALC_EXP_LOOP_and_svs_st_4;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0;
      COMPUTE_BATCH_LOOP_asn_2_itm_5 <= COMPUTE_BATCH_LOOP_asn_2_itm_4;
      CALC_EXP_LOOP_and_svs_st_4 <= CALC_EXP_LOOP_and_svs_st_3;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0;
      COMPUTE_BATCH_LOOP_asn_2_itm_4 <= exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_3;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_3 <= exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_2;
      CALC_SOFTMAX_LOOP_asn_itm_3 <= CALC_SOFTMAX_LOOP_asn_itm_2;
      CALC_EXP_LOOP_and_svs_st_2 <= CALC_EXP_LOOP_and_svs_st_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_2 <= exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_1;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_1 <= ~ COMPUTE_BATCH_LOOP_acc_itm_32_1;
      CALC_SOFTMAX_LOOP_asn_itm_1 <= exitL_exit_CALC_SOFTMAX_LOOP_sva;
      COMPUTE_BATCH_LOOP_stage_0 <= ~((~(COMPUTE_BATCH_LOOP_stage_0 & (COMPUTE_BATCH_LOOP_acc_itm_32_1
          | (~ exitL_exit_CALC_SOFTMAX_LOOP_sva)))) & (fsm_output[1]));
      exitL_exit_CALC_SOFTMAX_LOOP_sva <= ~((lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1_1
          | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0_1) & (fsm_output[1]));
      COMPUTE_BATCH_LOOP_stage_0_2 <= COMPUTE_BATCH_LOOP_stage_0 & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_3 <= COMPUTE_BATCH_LOOP_stage_0_2 & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_4 <= COMPUTE_BATCH_LOOP_stage_0_3 & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_5 <= COMPUTE_BATCH_LOOP_stage_0_4 & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_6 <= COMPUTE_BATCH_LOOP_stage_0_5 & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_7 <= COMPUTE_BATCH_LOOP_stage_0_6 & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_8 <= COMPUTE_BATCH_LOOP_stage_0_7 & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_9 <= COMPUTE_BATCH_LOOP_stage_0_8 & (fsm_output[1]);
      COMPUTE_BATCH_LOOP_stage_0_10 <= COMPUTE_BATCH_LOOP_stage_0_9 & (fsm_output[1]);
      ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_itm_1
          <= ~((SUM_EXP_LOOP_acc_1_tmp!=74'b00000000000000000000000000000000000000000000000000000000000000000000000000));
      CALC_SOFTMAX_LOOP_and_10_itm_5 <= CALC_SOFTMAX_LOOP_and_10_itm_4;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_4 <= CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_3;
      exit_COMPUTE_BATCH_LOOP_sva_1_3 <= exit_COMPUTE_BATCH_LOOP_sva_1_2;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_7 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_6;
      CALC_EXP_LOOP_and_svs_st_1 <= MUX_s_1_2_2(and_76_cse, (CALC_SOFTMAX_LOOP_acc_1_tmp[7]),
          and_dcpl_77);
      CALC_EXP_LOOP_and_svs_st_3 <= CALC_EXP_LOOP_and_svs_st_2;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1_mx0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0_mx0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_1 <= (~ COMPUTE_BATCH_LOOP_acc_itm_32_1)
          & exitL_exit_CALC_SOFTMAX_LOOP_sva;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_7 <= exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_6;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_6 <= exit_COMPUTE_BATCH_LOOP_sva_1_st_5;
      CALC_SOFTMAX_LOOP_asn_itm_2 <= CALC_SOFTMAX_LOOP_asn_itm_1;
      CALC_SOFTMAX_LOOP_asn_itm_6 <= CALC_SOFTMAX_LOOP_asn_itm_5;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_6 <= CALC_EXP_LOOP_and_svs_st_5;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_0;
      exit_COMPUTE_BATCH_LOOP_lpi_1_dfm_st_6 <= COMPUTE_BATCH_LOOP_asn_2_itm_5;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_5 <= exit_COMPUTE_BATCH_LOOP_sva_1_st_4;
      CALC_SOFTMAX_LOOP_asn_itm_5 <= CALC_SOFTMAX_LOOP_asn_itm_4;
      CALC_SOFTMAX_LOOP_and_10_itm_4 <= CALC_SOFTMAX_LOOP_and_10_itm_3;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_3 <= CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_2;
      exit_COMPUTE_BATCH_LOOP_sva_1_2 <= exit_COMPUTE_BATCH_LOOP_sva_1_st_1;
      exit_COMPUTE_BATCH_LOOP_sva_1_st_4 <= exit_COMPUTE_BATCH_LOOP_sva_1_3;
      CALC_SOFTMAX_LOOP_asn_itm_4 <= CALC_SOFTMAX_LOOP_asn_itm_3;
      CALC_SOFTMAX_LOOP_and_10_itm_3 <= CALC_SOFTMAX_LOOP_and_10_itm_2;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_2 <= CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_1;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_1 <= CALC_SOFTMAX_LOOP_or_tmp_1;
      CALC_SOFTMAX_LOOP_and_10_itm_2 <= CALC_SOFTMAX_LOOP_and_10_itm_1;
      CALC_SOFTMAX_LOOP_and_10_itm_1 <= CALC_SOFTMAX_LOOP_and_5_ssc_1;
    end
  end
  always @(posedge clk) begin
    if ( ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_and_cse
        ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1
          <= MUX_v_94_2_2(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_or_nl,
          ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1,
          or_8_nl);
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1
          <= ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_mx1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0 <= 1'b0;
    end
    else if ( ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_and_cse
        ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_0_1;
    end
  end
  always @(posedge clk) begin
    if ( ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_and_cse ) begin
      ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm <= nl_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm[7:0];
      ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_slc_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_9_0_itm
          <= ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[9:0];
      ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm
          <= nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm[10:0];
    end
  end
  assign or_nl = exit_COMPUTE_BATCH_LOOP_sva_1_3 | (~ CALC_SOFTMAX_LOOP_asn_itm_3);
  assign nl_COMPUTE_BATCH_LOOP_acc_1_nl = COMPUTE_BATCH_LOOP_b_sva + 32'b00000000000000000000000000000001;
  assign COMPUTE_BATCH_LOOP_acc_1_nl = nl_COMPUTE_BATCH_LOOP_acc_1_nl[31:0];
  assign COMPUTE_BATCH_LOOP_b_and_nl = (exitL_exit_CALC_SOFTMAX_LOOP_sva | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_4_1)
      | (~ (CALC_SOFTMAX_LOOP_acc_1_tmp[7]))) & (fsm_output[1]);
  assign COMPUTE_BATCH_LOOP_b_mux_nl = MUX_v_32_2_2(COMPUTE_BATCH_LOOP_acc_1_nl,
      COMPUTE_BATCH_LOOP_b_sva, COMPUTE_BATCH_LOOP_b_and_nl);
  assign CALC_SOFTMAX_LOOP_and_14_nl = (~ CALC_SOFTMAX_LOOP_equal_tmp_2) & or_14_tmp;
  assign CALC_SOFTMAX_LOOP_and_15_nl = CALC_SOFTMAX_LOOP_equal_tmp_2 & or_14_tmp;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_or_nl
      = MUX_v_94_2_2(operator_94_21_false_AC_TRN_AC_WRAP_rshift_itm, 94'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
      ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_itm_1);
  assign or_8_nl = (~ COMPUTE_BATCH_LOOP_stage_0_6) | COMPUTE_BATCH_LOOP_asn_2_itm_5
      | (~ CALC_SOFTMAX_LOOP_and_10_itm_5);
  assign nl_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm  =
      ({1'b1 , (~ libraries_leading_sign_74_0_cfd8a2a1b60025d53198d215150438e7bf24_1)})
      + 8'b00110111;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl
      = MUX_v_10_8_2(10'b1111111101, 10'b1100011001, 10'b1001100100, 10'b0111010000,
      10'b0101010100, 10'b0011101011, 10'b0010010001, 10'b0001000100, operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm[72:70]);
  assign nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_itm
      = conv_s2u_9_11(ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:10])
      + ({1'b1 , ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl});

  function automatic [73:0] MUX1HOT_v_74_3_2;
    input [73:0] input_2;
    input [73:0] input_1;
    input [73:0] input_0;
    input [2:0] sel;
    reg [73:0] result;
  begin
    result = input_0 & {74{sel[0]}};
    result = result | ( input_1 & {74{sel[1]}});
    result = result | ( input_2 & {74{sel[2]}});
    MUX1HOT_v_74_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_8_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [9:0] input_2;
    input [9:0] input_3;
    input [9:0] input_4;
    input [9:0] input_5;
    input [9:0] input_6;
    input [9:0] input_7;
    input [2:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_10_8_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_4_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [1:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_3_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_4_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [4:0] input_2;
    input [4:0] input_3;
    input [1:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_5_4_2 = result;
  end
  endfunction


  function automatic [73:0] MUX_v_74_2_2;
    input [73:0] input_0;
    input [73:0] input_1;
    input [0:0] sel;
    reg [73:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_74_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_4_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [6:0] input_2;
    input [6:0] input_3;
    input [1:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_7_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_8_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2 = result;
  end
  endfunction


  function automatic [93:0] MUX_v_94_2_2;
    input [93:0] input_0;
    input [93:0] input_1;
    input [0:0] sel;
    reg [93:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_94_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [18:0] readslicef_47_19_28;
    input [46:0] vector;
    reg [46:0] tmp;
  begin
    tmp = vector >> 28;
    readslicef_47_19_28 = tmp[18:0];
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input [0:0] vector;
  begin
    signext_7_1= {{6{vector[0]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_s2u_9_11 = {{2{vector[8]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_11 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [18:0] conv_u2u_19_19 ;
    input [18:0]  vector ;
  begin
    conv_u2u_19_19 = vector;
  end
  endfunction


  function automatic [32:0] conv_u2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_33 = {1'b0, vector};
  end
  endfunction


  function automatic [73:0] conv_u2u_67_74 ;
    input [66:0]  vector ;
  begin
    conv_u2u_67_74 = {{7{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input (
  clk, rst, conf_info, dma_read_ctrl_val, dma_read_ctrl_rdy, dma_read_ctrl_msg, dma_read_chnl_val,
      dma_read_chnl_rdy, dma_read_chnl_msg, done, input_ready_req_req, input_ready_ack_ack,
      plm_in_cns_req_vz, plm_in_cns_rls_lz, plm_in_cnsi_d_d, plm_in_cnsi_wadr_d,
      plm_in_cnsi_we_d_pff
);
  input clk;
  input rst;
  input [31:0] conf_info;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  input done;
  output input_ready_req_req;
  input input_ready_ack_ack;
  input plm_in_cns_req_vz;
  output plm_in_cns_rls_lz;
  output [31:0] plm_in_cnsi_d_d;
  output [6:0] plm_in_cnsi_wadr_d;
  output plm_in_cnsi_we_d_pff;


  // Interconnect Declarations
  wire load_input_wen;
  wire load_input_wten;
  wire dma_read_ctrl_Push_mioi_wen_comp;
  wire dma_read_chnl_Pop_mioi_wen_comp;
  wire [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt;
  wire input_ready_req_mioi_wen_comp;
  wire plm_in_cns_req_obj_wen_comp;
  wire [2:0] fsm_output;
  wire [7:0] LOAD_DATA_INNER_LOOP_acc_1_tmp;
  wire [8:0] nl_LOAD_DATA_INNER_LOOP_acc_1_tmp;
  reg LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_7_1_itm_1;
  reg exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_1;
  reg LOAD_BATCH_LOOP_stage_0_2;
  reg LOAD_BATCH_LOOP_stage_0;
  reg exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2;
  reg LOAD_BATCH_LOOP_stage_0_3;
  reg LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_7_1_itm_2;
  reg reg_dma_read_ctrl_Push_mioi_oswt_cse;
  reg reg_dma_read_chnl_Pop_mioi_oswt_cse;
  reg reg_input_ready_req_mioi_oswt_cse;
  reg reg_plm_in_cns_rls_obj_iswt0_cse;
  wire or_7_cse;
  wire and_cse;
  wire plm_in_cnsi_we_d_iff;
  wire and_11_rmff;
  wire and_15_rmff;
  wire and_17_rmff;
  reg [6:0] LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_6_0_itm_1;
  reg [24:0] offset_31_7_sva;
  reg [31:0] config_batch_sva;
  reg [31:0] LOAD_BATCH_LOOP_b_sva;
  wire [6:0] LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_6_0_itm_1_mx0;
  reg [6:0] LOAD_DATA_INNER_LOOP_i_7_0_sva_1_6_0;
  wire LOAD_BATCH_LOOP_acc_itm_32_1;

  wire[24:0] offset_mux_nl;
  wire[24:0] LOAD_BATCH_LOOP_acc_1_nl;
  wire[25:0] nl_LOAD_BATCH_LOOP_acc_1_nl;
  wire[0:0] offset_and_nl;
  wire[31:0] LOAD_BATCH_LOOP_b_mux_nl;
  wire[31:0] LOAD_BATCH_LOOP_acc_2_nl;
  wire[32:0] nl_LOAD_BATCH_LOOP_acc_2_nl;
  wire[0:0] LOAD_BATCH_LOOP_b_and_nl;
  wire[32:0] LOAD_BATCH_LOOP_acc_nl;
  wire[33:0] nl_LOAD_BATCH_LOOP_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input;
  assign nl_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input
      = {offset_31_7_sva , 7'b0000000};
  wire [0:0] nl_softmax_load_input_load_input_plm_in_cnsi_1_inst_plm_in_cnsi_iswt0_pff;
  assign nl_softmax_load_input_load_input_plm_in_cnsi_1_inst_plm_in_cnsi_iswt0_pff
      = and_cse & (fsm_output[1]);
  wire [0:0] nl_softmax_load_input_load_input_plm_in_cnsi_1_inst_load_input_wten_pff;
  assign nl_softmax_load_input_load_input_plm_in_cnsi_1_inst_load_input_wten_pff
      = ~ load_input_wen;
  wire [0:0] nl_softmax_load_input_load_input_load_input_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  assign nl_softmax_load_input_load_input_load_input_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0
      = ~ done;
  wire [0:0] nl_softmax_load_input_load_input_load_input_fsm_inst_LOAD_BATCH_LOOP_C_0_tr0;
  assign nl_softmax_load_input_load_input_load_input_fsm_inst_LOAD_BATCH_LOOP_C_0_tr0
      = LOAD_BATCH_LOOP_stage_0_2 | LOAD_BATCH_LOOP_stage_0_3 | LOAD_BATCH_LOOP_stage_0;
  esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi softmax_load_input_load_input_dma_read_ctrl_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_ctrl_val(dma_read_ctrl_val),
      .dma_read_ctrl_rdy(dma_read_ctrl_rdy),
      .dma_read_ctrl_msg(dma_read_ctrl_msg),
      .load_input_wen(load_input_wen),
      .dma_read_ctrl_Push_mioi_oswt(reg_dma_read_ctrl_Push_mioi_oswt_cse),
      .dma_read_ctrl_Push_mioi_wen_comp(dma_read_ctrl_Push_mioi_wen_comp),
      .dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input(nl_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input[31:0]),
      .dma_read_ctrl_Push_mioi_oswt_pff(and_11_rmff)
    );
  esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi softmax_load_input_load_input_dma_read_chnl_Pop_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_chnl_val(dma_read_chnl_val),
      .dma_read_chnl_rdy(dma_read_chnl_rdy),
      .dma_read_chnl_msg(dma_read_chnl_msg),
      .load_input_wen(load_input_wen),
      .dma_read_chnl_Pop_mioi_oswt(reg_dma_read_chnl_Pop_mioi_oswt_cse),
      .dma_read_chnl_Pop_mioi_wen_comp(dma_read_chnl_Pop_mioi_wen_comp),
      .dma_read_chnl_Pop_mioi_return_rsc_z_mxwt(dma_read_chnl_Pop_mioi_return_rsc_z_mxwt),
      .dma_read_chnl_Pop_mioi_oswt_pff(and_15_rmff)
    );
  esp_acc_softmax_softmax_load_input_load_input_input_ready_req_mioi softmax_load_input_load_input_input_ready_req_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .input_ready_req_req(input_ready_req_req),
      .input_ready_ack_ack(input_ready_ack_ack),
      .load_input_wen(load_input_wen),
      .input_ready_req_mioi_oswt(reg_input_ready_req_mioi_oswt_cse),
      .input_ready_req_mioi_wen_comp(input_ready_req_mioi_wen_comp),
      .input_ready_req_mioi_oswt_pff(and_17_rmff)
    );
  esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi_1 softmax_load_input_load_input_plm_in_cnsi_1_inst
      (
      .plm_in_cnsi_we_d_pff(plm_in_cnsi_we_d_iff),
      .plm_in_cnsi_iswt0_pff(nl_softmax_load_input_load_input_plm_in_cnsi_1_inst_plm_in_cnsi_iswt0_pff[0:0]),
      .load_input_wten_pff(nl_softmax_load_input_load_input_plm_in_cnsi_1_inst_load_input_wten_pff[0:0])
    );
  esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_rls_obj softmax_load_input_load_input_plm_in_cns_rls_obj_inst
      (
      .plm_in_cns_rls_lz(plm_in_cns_rls_lz),
      .load_input_wten(load_input_wten),
      .plm_in_cns_rls_obj_iswt0(reg_plm_in_cns_rls_obj_iswt0_cse)
    );
  esp_acc_softmax_softmax_load_input_load_input_plm_in_cns_req_obj softmax_load_input_load_input_plm_in_cns_req_obj_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_req_vz(plm_in_cns_req_vz),
      .load_input_wen(load_input_wen),
      .plm_in_cns_req_obj_oswt(reg_dma_read_ctrl_Push_mioi_oswt_cse),
      .plm_in_cns_req_obj_wen_comp(plm_in_cns_req_obj_wen_comp)
    );
  esp_acc_softmax_softmax_load_input_load_input_staller softmax_load_input_load_input_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .load_input_wen(load_input_wen),
      .load_input_wten(load_input_wten),
      .dma_read_ctrl_Push_mioi_wen_comp(dma_read_ctrl_Push_mioi_wen_comp),
      .dma_read_chnl_Pop_mioi_wen_comp(dma_read_chnl_Pop_mioi_wen_comp),
      .input_ready_req_mioi_wen_comp(input_ready_req_mioi_wen_comp),
      .plm_in_cns_req_obj_wen_comp(plm_in_cns_req_obj_wen_comp)
    );
  esp_acc_softmax_softmax_load_input_load_input_load_input_fsm softmax_load_input_load_input_load_input_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .load_input_wen(load_input_wen),
      .fsm_output(fsm_output),
      .WAIT_FOR_CONFIG_LOOP_C_0_tr0(nl_softmax_load_input_load_input_load_input_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0[0:0]),
      .LOAD_BATCH_LOOP_C_0_tr0(nl_softmax_load_input_load_input_load_input_fsm_inst_LOAD_BATCH_LOOP_C_0_tr0[0:0])
    );
  assign and_11_rmff = LOAD_BATCH_LOOP_acc_itm_32_1 & LOAD_BATCH_LOOP_stage_0 & LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_7_1_itm_1
      & (fsm_output[1]);
  assign and_15_rmff = or_7_cse & LOAD_BATCH_LOOP_stage_0 & (fsm_output[1]);
  assign and_17_rmff = LOAD_BATCH_LOOP_stage_0_3 & LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_7_1_itm_2
      & (~ exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2) & (fsm_output[1]);
  assign and_cse = LOAD_BATCH_LOOP_stage_0_2 & (~ exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_1);
  assign or_7_cse = LOAD_BATCH_LOOP_acc_itm_32_1 | (~ LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_7_1_itm_1);
  assign LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_6_0_itm_1_mx0 = MUX_v_7_2_2(LOAD_DATA_INNER_LOOP_i_7_0_sva_1_6_0,
      (signext_7_1(~ LOAD_BATCH_LOOP_acc_itm_32_1)), LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_7_1_itm_1);
  assign nl_LOAD_DATA_INNER_LOOP_acc_1_tmp = conv_u2u_7_8(LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_6_0_itm_1_mx0)
      + 8'b00000001;
  assign LOAD_DATA_INNER_LOOP_acc_1_tmp = nl_LOAD_DATA_INNER_LOOP_acc_1_tmp[7:0];
  assign nl_LOAD_BATCH_LOOP_acc_nl = ({1'b1 , LOAD_BATCH_LOOP_b_sva}) + conv_u2u_32_33(~
      config_batch_sva) + 33'b000000000000000000000000000000001;
  assign LOAD_BATCH_LOOP_acc_nl = nl_LOAD_BATCH_LOOP_acc_nl[32:0];
  assign LOAD_BATCH_LOOP_acc_itm_32_1 = readslicef_33_1_32(LOAD_BATCH_LOOP_acc_nl);
  assign plm_in_cnsi_d_d = dma_read_chnl_Pop_mioi_return_rsc_z_mxwt;
  assign plm_in_cnsi_wadr_d = LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_6_0_itm_1;
  assign plm_in_cnsi_we_d_pff = plm_in_cnsi_we_d_iff;
  always @(posedge clk) begin
    if ( load_input_wen ) begin
      LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_6_0_itm_1 <= LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_6_0_itm_1_mx0;
      offset_31_7_sva <= MUX_v_25_2_2(25'b0000000000000000000000000, offset_mux_nl,
          (fsm_output[1]));
      LOAD_BATCH_LOOP_b_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          LOAD_BATCH_LOOP_b_mux_nl, (fsm_output[1]));
      config_batch_sva <= MUX_v_32_2_2(conf_info, config_batch_sva, fsm_output[1]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_dma_read_ctrl_Push_mioi_oswt_cse <= 1'b0;
      reg_dma_read_chnl_Pop_mioi_oswt_cse <= 1'b0;
      reg_input_ready_req_mioi_oswt_cse <= 1'b0;
      reg_plm_in_cns_rls_obj_iswt0_cse <= 1'b0;
      LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_7_1_itm_2 <= 1'b0;
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2 <= 1'b0;
      LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_7_1_itm_1 <= 1'b0;
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_1 <= 1'b0;
      LOAD_BATCH_LOOP_stage_0 <= 1'b0;
      LOAD_DATA_INNER_LOOP_i_7_0_sva_1_6_0 <= 7'b0000000;
      LOAD_BATCH_LOOP_stage_0_2 <= 1'b0;
      LOAD_BATCH_LOOP_stage_0_3 <= 1'b0;
    end
    else if ( load_input_wen ) begin
      reg_dma_read_ctrl_Push_mioi_oswt_cse <= and_11_rmff;
      reg_dma_read_chnl_Pop_mioi_oswt_cse <= and_15_rmff;
      reg_input_ready_req_mioi_oswt_cse <= and_17_rmff;
      reg_plm_in_cns_rls_obj_iswt0_cse <= and_cse & LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_7_1_itm_1
          & (fsm_output[1]);
      LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_7_1_itm_2 <= LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_7_1_itm_1;
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_2 <= exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_1;
      LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_7_1_itm_1 <= (LOAD_DATA_INNER_LOOP_acc_1_tmp[7])
          | (~ (fsm_output[1]));
      exit_LOAD_BATCH_LOOP_lpi_1_dfm_st_1 <= (~ LOAD_BATCH_LOOP_acc_itm_32_1) & LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_7_1_itm_1;
      LOAD_BATCH_LOOP_stage_0 <= ~((~(LOAD_BATCH_LOOP_stage_0 & or_7_cse)) & (fsm_output[1]));
      LOAD_DATA_INNER_LOOP_i_7_0_sva_1_6_0 <= LOAD_DATA_INNER_LOOP_acc_1_tmp[6:0];
      LOAD_BATCH_LOOP_stage_0_2 <= LOAD_BATCH_LOOP_stage_0 & (fsm_output[1]);
      LOAD_BATCH_LOOP_stage_0_3 <= LOAD_BATCH_LOOP_stage_0_2 & (fsm_output[1]);
    end
  end
  assign nl_LOAD_BATCH_LOOP_acc_1_nl = offset_31_7_sva + 25'b0000000000000000000000001;
  assign LOAD_BATCH_LOOP_acc_1_nl = nl_LOAD_BATCH_LOOP_acc_1_nl[24:0];
  assign offset_and_nl = LOAD_DATA_INNER_LOOP_i_slc_LOAD_DATA_INNER_LOOP_i_7_0_7_1_itm_1
      & (fsm_output[1]);
  assign offset_mux_nl = MUX_v_25_2_2(offset_31_7_sva, LOAD_BATCH_LOOP_acc_1_nl,
      offset_and_nl);
  assign nl_LOAD_BATCH_LOOP_acc_2_nl = LOAD_BATCH_LOOP_b_sva + 32'b00000000000000000000000000000001;
  assign LOAD_BATCH_LOOP_acc_2_nl = nl_LOAD_BATCH_LOOP_acc_2_nl[31:0];
  assign LOAD_BATCH_LOOP_b_and_nl = (LOAD_DATA_INNER_LOOP_acc_1_tmp[7]) & (fsm_output[1]);
  assign LOAD_BATCH_LOOP_b_mux_nl = MUX_v_32_2_2(LOAD_BATCH_LOOP_b_sva, LOAD_BATCH_LOOP_acc_2_nl,
      LOAD_BATCH_LOOP_b_and_nl);

  function automatic [24:0] MUX_v_25_2_2;
    input [24:0] input_0;
    input [24:0] input_1;
    input [0:0] sel;
    reg [24:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_25_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input [0:0] vector;
  begin
    signext_7_1= {{6{vector[0]}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [32:0] conv_u2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_33 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output (
  clk, rst, conf_info, acc_done, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg,
      dma_write_chnl_val, dma_write_chnl_rdy, dma_write_chnl_msg, done, output_ready_req_req,
      output_ready_ack_ack, plm_out_cns_radr, plm_out_cns_q, plm_out_cns_req_vz,
      plm_out_cns_rls_lz
);
  input clk;
  input rst;
  input [31:0] conf_info;
  output acc_done;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;
  input done;
  input output_ready_req_req;
  output output_ready_ack_ack;
  output [6:0] plm_out_cns_radr;
  input [31:0] plm_out_cns_q;
  input plm_out_cns_req_vz;
  output plm_out_cns_rls_lz;


  // Interconnect Declarations
  wire [31:0] plm_out_cnsi_q_d;
  wire [6:0] plm_out_cnsi_radr_d;
  wire plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_softmax_store_output_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_40_7_32_128_128_32_1_gen
      plm_out_cnsi (
      .q(plm_out_cns_q),
      .radr(plm_out_cns_radr),
      .q_d(plm_out_cnsi_q_d),
      .radr_d(plm_out_cnsi_radr_d),
      .readA_r_ram_ir_internal_RMASK_B_d(plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_softmax_softmax_store_output_store_output softmax_store_output_store_output_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .acc_done(acc_done),
      .dma_write_ctrl_val(dma_write_ctrl_val),
      .dma_write_ctrl_rdy(dma_write_ctrl_rdy),
      .dma_write_ctrl_msg(dma_write_ctrl_msg),
      .dma_write_chnl_val(dma_write_chnl_val),
      .dma_write_chnl_rdy(dma_write_chnl_rdy),
      .dma_write_chnl_msg(dma_write_chnl_msg),
      .done(done),
      .output_ready_req_req(output_ready_req_req),
      .output_ready_ack_ack(output_ready_ack_ack),
      .plm_out_cns_req_vz(plm_out_cns_req_vz),
      .plm_out_cns_rls_lz(plm_out_cns_rls_lz),
      .plm_out_cnsi_q_d(plm_out_cnsi_q_d),
      .plm_out_cnsi_radr_d(plm_out_cnsi_radr_d),
      .plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d(plm_out_cnsi_readA_r_ram_ir_internal_RMASK_B_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel (
  clk, rst, conf_info, done, input_ready_req_req, input_ready_ack_ack, output_ready_req_req,
      output_ready_ack_ack, plm_in_cns_radr, plm_in_cns_q, plm_in_cns_req_vz, plm_in_cns_rls_lz,
      plm_out_cns_wadr, plm_out_cns_d, plm_out_cns_we, plm_out_cns_req_vz, plm_out_cns_rls_lz
);
  input clk;
  input rst;
  input [31:0] conf_info;
  input done;
  input input_ready_req_req;
  output input_ready_ack_ack;
  output output_ready_req_req;
  input output_ready_ack_ack;
  output [6:0] plm_in_cns_radr;
  input [31:0] plm_in_cns_q;
  input plm_in_cns_req_vz;
  output plm_in_cns_rls_lz;
  output [6:0] plm_out_cns_wadr;
  output [31:0] plm_out_cns_d;
  output plm_out_cns_we;
  input plm_out_cns_req_vz;
  output plm_out_cns_rls_lz;


  // Interconnect Declarations
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] plm_in_cnsi_q_d;
  wire [6:0] plm_in_cnsi_radr_d;
  wire plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d;
  wire [31:0] plm_out_cnsi_d_d;
  wire [6:0] plm_out_cnsi_wadr_d;
  wire [93:0] CALC_SOFTMAX_LOOP_mul_cmp_b;
  wire [94:0] CALC_SOFTMAX_LOOP_mul_cmp_z;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_clken;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_q;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_radr;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_we;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_d;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wadr;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d_iff;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff;
  wire plm_out_cnsi_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_mgc_mul_pipe #(.width_a(32'sd67),
  .signd_a(32'sd0),
  .width_b(32'sd94),
  .signd_b(32'sd0),
  .width_z(32'sd95),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) CALC_SOFTMAX_LOOP_mul_cmp (
      .a(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d),
      .b(CALC_SOFTMAX_LOOP_mul_cmp_b),
      .clk(clk),
      .en(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(CALC_SOFTMAX_LOOP_mul_cmp_z)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd7),
  .data_width(32'sd67),
  .depth(32'sd128),
  .latency(32'sd1)) ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_comp
      (
      .clk(clk),
      .clken(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_clken),
      .d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_d),
      .q(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_q),
      .radr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_radr),
      .wadr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wadr),
      .we(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_we)
    );
  esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_17_7_67_128_128_67_1_gen
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci
      (
      .clken(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_clken),
      .q(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_q),
      .radr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_radr),
      .we(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_we),
      .d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_d),
      .wadr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wadr),
      .clken_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d),
      .d_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d),
      .q_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d),
      .radr_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d_iff),
      .wadr_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d_iff),
      .we_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_34_7_32_128_128_32_1_gen
      plm_in_cnsi (
      .q(plm_in_cns_q),
      .radr(plm_in_cns_radr),
      .q_d(plm_in_cnsi_q_d),
      .radr_d(plm_in_cnsi_radr_d),
      .readA_r_ram_ir_internal_RMASK_B_d(plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_35_7_32_128_128_32_1_gen
      plm_out_cnsi (
      .we(plm_out_cns_we),
      .d(plm_out_cns_d),
      .wadr(plm_out_cns_wadr),
      .d_d(plm_out_cnsi_d_d),
      .wadr_d(plm_out_cnsi_wadr_d),
      .we_d(plm_out_cnsi_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(plm_out_cnsi_we_d_iff)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel softmax_compute_kernel_compute_kernel_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .done(done),
      .input_ready_req_req(input_ready_req_req),
      .input_ready_ack_ack(input_ready_ack_ack),
      .output_ready_req_req(output_ready_req_req),
      .output_ready_ack_ack(output_ready_ack_ack),
      .plm_in_cns_req_vz(plm_in_cns_req_vz),
      .plm_in_cns_rls_lz(plm_in_cns_rls_lz),
      .plm_out_cns_req_vz(plm_out_cns_req_vz),
      .plm_out_cns_rls_lz(plm_out_cns_rls_lz),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .plm_in_cnsi_q_d(plm_in_cnsi_q_d),
      .plm_in_cnsi_radr_d(plm_in_cnsi_radr_d),
      .plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d(plm_in_cnsi_readA_r_ram_ir_internal_RMASK_B_d),
      .plm_out_cnsi_d_d(plm_out_cnsi_d_d),
      .plm_out_cnsi_wadr_d(plm_out_cnsi_wadr_d),
      .CALC_SOFTMAX_LOOP_mul_cmp_b(CALC_SOFTMAX_LOOP_mul_cmp_b),
      .CALC_SOFTMAX_LOOP_mul_cmp_z(CALC_SOFTMAX_LOOP_mul_cmp_z),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d_pff(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d_iff),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff),
      .plm_out_cnsi_we_d_pff(plm_out_cnsi_we_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input (
  clk, rst, conf_info, dma_read_ctrl_val, dma_read_ctrl_rdy, dma_read_ctrl_msg, dma_read_chnl_val,
      dma_read_chnl_rdy, dma_read_chnl_msg, done, input_ready_req_req, input_ready_ack_ack,
      plm_in_cns_wadr, plm_in_cns_d, plm_in_cns_we, plm_in_cns_req_vz, plm_in_cns_rls_lz
);
  input clk;
  input rst;
  input [31:0] conf_info;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  input done;
  output input_ready_req_req;
  input input_ready_ack_ack;
  output [6:0] plm_in_cns_wadr;
  output [31:0] plm_in_cns_d;
  output plm_in_cns_we;
  input plm_in_cns_req_vz;
  output plm_in_cns_rls_lz;


  // Interconnect Declarations
  wire [31:0] plm_in_cnsi_d_d;
  wire [6:0] plm_in_cnsi_wadr_d;
  wire plm_in_cnsi_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_softmax_load_input_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_33_7_32_128_128_32_1_gen
      plm_in_cnsi (
      .we(plm_in_cns_we),
      .d(plm_in_cns_d),
      .wadr(plm_in_cns_wadr),
      .d_d(plm_in_cnsi_d_d),
      .wadr_d(plm_in_cnsi_wadr_d),
      .we_d(plm_in_cnsi_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(plm_in_cnsi_we_d_iff)
    );
  esp_acc_softmax_softmax_load_input_load_input softmax_load_input_load_input_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .dma_read_ctrl_val(dma_read_ctrl_val),
      .dma_read_ctrl_rdy(dma_read_ctrl_rdy),
      .dma_read_ctrl_msg(dma_read_ctrl_msg),
      .dma_read_chnl_val(dma_read_chnl_val),
      .dma_read_chnl_rdy(dma_read_chnl_rdy),
      .dma_read_chnl_msg(dma_read_chnl_msg),
      .done(done),
      .input_ready_req_req(input_ready_req_req),
      .input_ready_ack_ack(input_ready_ack_ack),
      .plm_in_cns_req_vz(plm_in_cns_req_vz),
      .plm_in_cns_rls_lz(plm_in_cns_rls_lz),
      .plm_in_cnsi_d_d(plm_in_cnsi_d_d),
      .plm_in_cnsi_wadr_d(plm_in_cnsi_wadr_d),
      .plm_in_cnsi_we_d_pff(plm_in_cnsi_we_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    softmax_basic_fx32_dma64
// ------------------------------------------------------------------


module softmax_basic_fx32_dma64 (
  clk, rst, conf_info, conf_done, acc_done, debug, dma_read_ctrl_val, dma_read_ctrl_rdy,
      dma_read_ctrl_msg, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg,
      dma_read_chnl_val, dma_read_chnl_rdy, dma_read_chnl_msg, dma_write_chnl_val,
      dma_write_chnl_rdy, dma_write_chnl_msg
);
  input clk;
  input rst;
  input [31:0] conf_info;
  input conf_done;
  output acc_done;
  output [31:0] debug;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;


  // Interconnect Declarations
  wire done;
  wire input_ready_req_req;
  wire input_ready_ack_ack;
  wire output_ready_req_req;
  wire output_ready_ack_ack;
  wire [6:0] plm_in_cns_wadr_nsoftmax_load_input_inst;
  wire [31:0] plm_in_cns_d_nsoftmax_load_input_inst;
  wire plm_in_cns_we_nsoftmax_load_input_inst;
  wire plm_in_cns_req_vz_nsoftmax_load_input_inst;
  wire [6:0] plm_in_cns_radr_nsoftmax_compute_kernel_inst;
  wire [31:0] plm_in_cns_q_nsoftmax_compute_kernel_inst;
  wire plm_in_cns_req_vz_nsoftmax_compute_kernel_inst;
  wire [6:0] plm_out_cns_wadr_nsoftmax_compute_kernel_inst;
  wire [31:0] plm_out_cns_d_nsoftmax_compute_kernel_inst;
  wire plm_out_cns_we_nsoftmax_compute_kernel_inst;
  wire plm_out_cns_req_vz_nsoftmax_compute_kernel_inst;
  wire plm_out_cns_we_nsoftmax_compute_kernel_inst_buz;
  wire [6:0] plm_out_cns_radr_nsoftmax_store_output_inst;
  wire [31:0] plm_out_cns_q_nsoftmax_store_output_inst;
  wire plm_out_cns_req_vz_nsoftmax_store_output_inst;
  wire plm_in_cns_rls_lz_nsoftmax_load_input_inst_bud;
  wire plm_in_cns_rls_lz_nsoftmax_compute_kernel_inst_bud;
  wire plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud;
  wire plm_out_cns_rls_lz_nsoftmax_compute_kernel_inst_bud;
  wire plm_out_cns_rls_lz_nsoftmax_store_output_inst_bud;
  wire plm_in_cns_R0;
  wire plm_in_cns_S1;
  wire plm_in_cns_R1;
  wire [31:0] plm_in_cns_d_shi0;
  wire [31:0] plm_in_cns_d_shi1;
  wire [31:0] plm_in_cns_q_sho0;
  wire [31:0] plm_in_cns_q_sho1;
  wire [6:0] plm_in_cns_radr_shi0;
  wire [6:0] plm_in_cns_radr_shi1;
  wire [6:0] plm_in_cns_wadr_shi0;
  wire [6:0] plm_in_cns_wadr_shi1;
  wire plm_in_cns_we_shi0;
  wire plm_in_cns_we_shi1;
  wire plm_out_cns_R0;
  wire plm_out_cns_S1;
  wire plm_out_cns_R1;
  wire [31:0] plm_out_cns_d_shi0;
  wire [31:0] plm_out_cns_d_shi1;
  wire [31:0] plm_out_cns_q_sho0;
  wire [31:0] plm_out_cns_q_sho1;
  wire [6:0] plm_out_cns_radr_shi0;
  wire [6:0] plm_out_cns_radr_shi1;
  wire [6:0] plm_out_cns_wadr_shi0;
  wire [6:0] plm_out_cns_wadr_shi1;
  wire plm_out_cns_we_shi0;
  wire plm_out_cns_we_shi1;
  wire plm_in_cns_S0_iff;
  wire plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_iff;
  wire plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud_iff;
  wire plm_out_cns_S0_iff;
  wire plm_in_cns_S0_dmo;
  wire plm_out_cns_S0_dmo;


  // Interconnect Declarations for Component Instantiations 
  BLOCK_1R1W_RBW #(.addr_width(32'sd7),
  .data_width(32'sd32),
  .depth(32'sd128),
  .latency(32'sd1)) plm_in_cns_comp (
      .clk(clk),
      .clken(1'b1),
      .d(plm_in_cns_d_shi0),
      .q(plm_in_cns_q_sho0),
      .radr(plm_in_cns_radr_shi0),
      .wadr(plm_in_cns_wadr_shi0),
      .we(plm_in_cns_we_shi0)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd7),
  .data_width(32'sd32),
  .depth(32'sd128),
  .latency(32'sd1)) plm_in_cns_comp_1 (
      .clk(clk),
      .clken(1'b1),
      .d(plm_in_cns_d_shi1),
      .q(plm_in_cns_q_sho1),
      .radr(plm_in_cns_radr_shi1),
      .wadr(plm_in_cns_wadr_shi1),
      .we(plm_in_cns_we_shi1)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd7),
  .data_width(32'sd32),
  .depth(32'sd128),
  .latency(32'sd1)) plm_out_cns_comp (
      .clk(clk),
      .clken(1'b1),
      .d(plm_out_cns_d_shi0),
      .q(plm_out_cns_q_sho0),
      .radr(plm_out_cns_radr_shi0),
      .wadr(plm_out_cns_wadr_shi0),
      .we(plm_out_cns_we_shi0)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd7),
  .data_width(32'sd32),
  .depth(32'sd128),
  .latency(32'sd1)) plm_out_cns_comp_1 (
      .clk(clk),
      .clken(1'b1),
      .d(plm_out_cns_d_shi1),
      .q(plm_out_cns_q_sho1),
      .radr(plm_out_cns_radr_shi1),
      .wadr(plm_out_cns_wadr_shi1),
      .we(plm_out_cns_we_shi1)
    );
  esp_acc_softmax_softmax_load_input softmax_load_input_inst (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .dma_read_ctrl_val(dma_read_ctrl_val),
      .dma_read_ctrl_rdy(dma_read_ctrl_rdy),
      .dma_read_ctrl_msg(dma_read_ctrl_msg),
      .dma_read_chnl_val(dma_read_chnl_val),
      .dma_read_chnl_rdy(dma_read_chnl_rdy),
      .dma_read_chnl_msg(dma_read_chnl_msg),
      .done(done),
      .input_ready_req_req(input_ready_req_req),
      .input_ready_ack_ack(input_ready_ack_ack),
      .plm_in_cns_wadr(plm_in_cns_wadr_nsoftmax_load_input_inst),
      .plm_in_cns_d(plm_in_cns_d_nsoftmax_load_input_inst),
      .plm_in_cns_we(plm_in_cns_we_nsoftmax_load_input_inst),
      .plm_in_cns_req_vz(plm_in_cns_req_vz_nsoftmax_load_input_inst),
      .plm_in_cns_rls_lz(plm_in_cns_rls_lz_nsoftmax_load_input_inst_bud)
    );
  esp_acc_softmax_softmax_compute_kernel softmax_compute_kernel_inst (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .done(done),
      .input_ready_req_req(input_ready_req_req),
      .input_ready_ack_ack(input_ready_ack_ack),
      .output_ready_req_req(output_ready_req_req),
      .output_ready_ack_ack(output_ready_ack_ack),
      .plm_in_cns_radr(plm_in_cns_radr_nsoftmax_compute_kernel_inst),
      .plm_in_cns_q(plm_in_cns_q_nsoftmax_compute_kernel_inst),
      .plm_in_cns_req_vz(plm_in_cns_req_vz_nsoftmax_compute_kernel_inst),
      .plm_in_cns_rls_lz(plm_in_cns_rls_lz_nsoftmax_compute_kernel_inst_bud),
      .plm_out_cns_wadr(plm_out_cns_wadr_nsoftmax_compute_kernel_inst),
      .plm_out_cns_d(plm_out_cns_d_nsoftmax_compute_kernel_inst),
      .plm_out_cns_we(plm_out_cns_we_nsoftmax_compute_kernel_inst),
      .plm_out_cns_req_vz(plm_out_cns_req_vz_nsoftmax_compute_kernel_inst),
      .plm_out_cns_rls_lz(plm_out_cns_rls_lz_nsoftmax_compute_kernel_inst_bud)
    );
  esp_acc_softmax_softmax_store_output softmax_store_output_inst (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .acc_done(acc_done),
      .dma_write_ctrl_val(dma_write_ctrl_val),
      .dma_write_ctrl_rdy(dma_write_ctrl_rdy),
      .dma_write_ctrl_msg(dma_write_ctrl_msg),
      .dma_write_chnl_val(dma_write_chnl_val),
      .dma_write_chnl_rdy(dma_write_chnl_rdy),
      .dma_write_chnl_msg(dma_write_chnl_msg),
      .done(done),
      .output_ready_req_req(output_ready_req_req),
      .output_ready_ack_ack(output_ready_ack_ack),
      .plm_out_cns_radr(plm_out_cns_radr_nsoftmax_store_output_inst),
      .plm_out_cns_q(plm_out_cns_q_nsoftmax_store_output_inst),
      .plm_out_cns_req_vz(plm_out_cns_req_vz_nsoftmax_store_output_inst),
      .plm_out_cns_rls_lz(plm_out_cns_rls_lz_nsoftmax_store_output_inst_bud)
    );
  esp_acc_softmax_unreg_hier unreg (
      .in_0(plm_in_cns_S0_iff),
      .out_0(plm_in_cns_R0)
    );
  esp_acc_softmax_unreg_hier unreg_1 (
      .in_0(plm_in_cns_S1),
      .out_0(plm_in_cns_R1)
    );
  esp_acc_softmax_unreg_hier unreg_2 (
      .in_0(plm_out_cns_S0_iff),
      .out_0(plm_out_cns_R0)
    );
  esp_acc_softmax_unreg_hier unreg_3 (
      .in_0(plm_out_cns_S1),
      .out_0(plm_out_cns_R1)
    );
  esp_acc_softmax_softmax_plm_in_cns_bctl softmax_plm_in_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_wadr_nsoftmax_load_input_inst(plm_in_cns_wadr_nsoftmax_load_input_inst),
      .plm_in_cns_d_nsoftmax_load_input_inst(plm_in_cns_d_nsoftmax_load_input_inst),
      .plm_in_cns_we_nsoftmax_load_input_inst(plm_in_cns_we_nsoftmax_load_input_inst),
      .plm_in_cns_req_vz_nsoftmax_load_input_inst(plm_in_cns_req_vz_nsoftmax_load_input_inst),
      .plm_in_cns_radr_nsoftmax_compute_kernel_inst(plm_in_cns_radr_nsoftmax_compute_kernel_inst),
      .plm_in_cns_q_nsoftmax_compute_kernel_inst(plm_in_cns_q_nsoftmax_compute_kernel_inst),
      .plm_in_cns_req_vz_nsoftmax_compute_kernel_inst(plm_in_cns_req_vz_nsoftmax_compute_kernel_inst),
      .plm_out_cns_we_nsoftmax_compute_kernel_inst_buz(plm_out_cns_we_nsoftmax_compute_kernel_inst_buz),
      .plm_in_cns_rls_lz_nsoftmax_load_input_inst_bud(plm_in_cns_rls_lz_nsoftmax_load_input_inst_bud),
      .plm_in_cns_rls_lz_nsoftmax_compute_kernel_inst_bud(plm_in_cns_rls_lz_nsoftmax_compute_kernel_inst_bud),
      .plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud(plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud),
      .plm_out_cns_rls_lz_nsoftmax_compute_kernel_inst_bud(1'b0),
      .plm_in_cns_S0(plm_in_cns_S0_dmo),
      .plm_in_cns_R0(plm_in_cns_R0),
      .plm_in_cns_S1(plm_in_cns_S1),
      .plm_in_cns_R1(plm_in_cns_R1),
      .plm_in_cns_d_shi0(plm_in_cns_d_shi0),
      .plm_in_cns_d_shi1(plm_in_cns_d_shi1),
      .plm_in_cns_q_sho0(plm_in_cns_q_sho0),
      .plm_in_cns_q_sho1(plm_in_cns_q_sho1),
      .plm_in_cns_radr_shi0(plm_in_cns_radr_shi0),
      .plm_in_cns_radr_shi1(plm_in_cns_radr_shi1),
      .plm_in_cns_wadr_shi0(plm_in_cns_wadr_shi0),
      .plm_in_cns_wadr_shi1(plm_in_cns_wadr_shi1),
      .plm_in_cns_we_shi0(plm_in_cns_we_shi0),
      .plm_in_cns_we_shi1(plm_in_cns_we_shi1),
      .plm_in_cns_S0_pff(plm_in_cns_S0_iff),
      .plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_pff(plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_iff),
      .plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud_pff(plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud_iff)
    );
  esp_acc_softmax_softmax_plm_out_cns_bctl softmax_plm_out_cns_bctl_inst (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_wadr_nsoftmax_compute_kernel_inst(plm_out_cns_wadr_nsoftmax_compute_kernel_inst),
      .plm_out_cns_d_nsoftmax_compute_kernel_inst(plm_out_cns_d_nsoftmax_compute_kernel_inst),
      .plm_out_cns_we_nsoftmax_compute_kernel_inst(plm_out_cns_we_nsoftmax_compute_kernel_inst),
      .plm_out_cns_req_vz_nsoftmax_compute_kernel_inst(plm_out_cns_req_vz_nsoftmax_compute_kernel_inst),
      .plm_out_cns_we_nsoftmax_compute_kernel_inst_buz(1'b0),
      .plm_out_cns_radr_nsoftmax_store_output_inst(plm_out_cns_radr_nsoftmax_store_output_inst),
      .plm_out_cns_q_nsoftmax_store_output_inst(plm_out_cns_q_nsoftmax_store_output_inst),
      .plm_out_cns_req_vz_nsoftmax_store_output_inst(plm_out_cns_req_vz_nsoftmax_store_output_inst),
      .plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud(plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud),
      .plm_out_cns_rls_lz_nsoftmax_compute_kernel_inst_bud(plm_out_cns_rls_lz_nsoftmax_compute_kernel_inst_bud),
      .plm_out_cns_rls_lz_nsoftmax_store_output_inst_bud(plm_out_cns_rls_lz_nsoftmax_store_output_inst_bud),
      .plm_out_cns_S0(plm_out_cns_S0_dmo),
      .plm_out_cns_R0(plm_out_cns_R0),
      .plm_out_cns_S1(plm_out_cns_S1),
      .plm_out_cns_R1(plm_out_cns_R1),
      .plm_out_cns_d_shi0(plm_out_cns_d_shi0),
      .plm_out_cns_d_shi1(plm_out_cns_d_shi1),
      .plm_out_cns_q_sho0(plm_out_cns_q_sho0),
      .plm_out_cns_q_sho1(plm_out_cns_q_sho1),
      .plm_out_cns_radr_shi0(plm_out_cns_radr_shi0),
      .plm_out_cns_radr_shi1(plm_out_cns_radr_shi1),
      .plm_out_cns_wadr_shi0(plm_out_cns_wadr_shi0),
      .plm_out_cns_wadr_shi1(plm_out_cns_wadr_shi1),
      .plm_out_cns_we_shi0(plm_out_cns_we_shi0),
      .plm_out_cns_we_shi1(plm_out_cns_we_shi1),
      .plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_pff(plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_iff),
      .plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud_pff(plm_out_cns_we_nsoftmax_compute_kernel_inst_buz_bud_iff),
      .plm_out_cns_S0_pff(plm_out_cns_S0_iff)
    );
  esp_acc_softmax_softmax_config_accelerator softmax_config_accelerator_inst (
      .clk(clk),
      .rst(rst),
      .conf_done(conf_done),
      .done(done)
    );
  assign debug = 32'b00000000000000000000000000000000;
endmodule



