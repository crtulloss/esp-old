
//------> ./softmax_Connections_OutBlockingless_dma_info_tcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_Connections_OutBlockingless_dma_info_tcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_Connections_OutBlockingless_dma_info_tcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Sun May  3 17:05:16 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core
    (
  this_val, this_rdy, this_msg, m_index_rsc_dat, m_length_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [66:0] this_msg;
  input [31:0] m_index_rsc_dat;
  input [31:0] m_length_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire [31:0] m_index_rsci_idat;
  wire [31:0] m_length_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [31:0] m_length_buf_lpi_1_dfm;
  reg [31:0] m_index_buf_lpi_1_dfm;
  wire and_dcpl;
  wire or_dcpl_2;
  reg LOAD_DATA_OUTER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire LOAD_DATA_OUTER_LOOP_LOAD_DATA_OUTER_LOOP_or_cse;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = LOAD_DATA_OUTER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd32)) m_index_rsci (
      .dat(m_index_rsc_dat),
      .idat(m_index_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd32)) m_length_rsci (
      .dat(m_length_rsc_dat),
      .idat(m_length_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd47),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 #(.rscid(32'sd56)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign this_msg = {3'b000 , m_length_buf_lpi_1_dfm , m_index_buf_lpi_1_dfm};
  assign LOAD_DATA_OUTER_LOOP_LOAD_DATA_OUTER_LOOP_or_cse = ccs_ccore_start_rsci_idat
      | and_dcpl;
  assign and_dcpl = LOAD_DATA_OUTER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_rdy);
  assign or_dcpl_2 = and_dcpl | (~ ccs_ccore_start_rsci_idat);
  assign this_val_mx0c1 = LOAD_DATA_OUTER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_val <= 1'b0;
    end
    else if ( LOAD_DATA_OUTER_LOOP_LOAD_DATA_OUTER_LOOP_or_cse | this_val_mx0c1 )
        begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      m_length_buf_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_length_buf_lpi_1_dfm <= m_length_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      m_index_buf_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~ or_dcpl_2 ) begin
      m_index_buf_lpi_1_dfm <= m_index_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      LOAD_DATA_OUTER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      LOAD_DATA_OUTER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= LOAD_DATA_OUTER_LOOP_LOAD_DATA_OUTER_LOOP_or_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module esp_acc_softmax_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_index_rsc_dat, m_length_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  input this_rdy;
  output [66:0] this_msg;
  input [31:0] m_index_rsc_dat;
  input [31:0] m_length_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_esp_acc_softmax_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core_inst (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_index_rsc_dat(m_index_rsc_dat),
      .m_length_rsc_dat(m_length_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_Connections_InBlockingless_sc_dt_sc_bvless_64greater_comma_Connections_SYN_PORTgreater_Pop_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./softmax_Connections_InBlockingless_sc_dt_sc_bvless_64greater_comma_Connections_SYN_PORTgreater_Pop_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_Connections_InBlockingless_sc_dt_sc_bvless_64greater_comma_Connections_SYN_PORTgreater_Pop_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_Connections_InBlockingless_sc_dt_sc_bvless_64greater_comma_Connections_SYN_PORTgreater_Pop.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Sun May  3 17:05:20 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_Connections_InBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Pop_core
// ------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_Connections_InBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Pop_core
    (
  this_val, this_rdy, this_msg, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [63:0] this_msg;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg LOAD_DATA_INNER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire LOAD_DATA_INNER_LOOP_LOAD_DATA_INNER_LOOP_or_cse;
  wire this_rdy_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [63:0] nl_return_rsci_d;
  assign nl_return_rsci_d = this_msg;
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = LOAD_DATA_INNER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_val;
  esp_acc_softmax_esp_acc_softmax_mgc_out_dreg_v2 #(.rscid(32'sd4),
  .width(32'sd64)) return_rsci (
      .d(nl_return_rsci_d[63:0]),
      .z(return_rsc_z)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd46),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 #(.rscid(32'sd55)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign LOAD_DATA_INNER_LOOP_LOAD_DATA_INNER_LOOP_or_cse = ccs_ccore_start_rsci_idat
      | (LOAD_DATA_INNER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_val));
  assign this_rdy_mx0c1 = LOAD_DATA_INNER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_val & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_rdy <= 1'b0;
    end
    else if ( LOAD_DATA_INNER_LOOP_LOAD_DATA_INNER_LOOP_or_cse | this_rdy_mx0c1 )
        begin
      this_rdy <= ~ this_rdy_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      LOAD_DATA_INNER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      LOAD_DATA_INNER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= LOAD_DATA_INNER_LOOP_LOAD_DATA_INNER_LOOP_or_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Pop
// ------------------------------------------------------------------


module esp_acc_softmax_Connections_InBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Pop (
  this_val, this_rdy, this_msg, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  input this_val;
  output this_rdy;
  input [63:0] this_msg;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_esp_acc_softmax_Connections_InBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Pop_core
      Connections_InBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Pop_core_inst (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_Connections_Combinationalless_boolcomma_Connections_SYN_PORTgreater_Pop_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./softmax_Connections_Combinationalless_boolcomma_Connections_SYN_PORTgreater_Pop_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_Connections_Combinationalless_boolcomma_Connections_SYN_PORTgreater_Pop_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_Connections_Combinationalless_boolcomma_Connections_SYN_PORTgreater_Pop.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Sun May  3 17:05:18 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_Connections_Combinational_bool_Connections_SYN_PORT_Pop_core
// ------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_Connections_Combinational_bool_Connections_SYN_PORT_Pop_core
    (
  this_val, this_rdy, this_msg, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input this_msg;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg input_ready_req_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire input_ready_req_input_ready_req_or_cse;
  wire this_rdy_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_return_rsci_d;
  assign nl_return_rsci_d = this_msg;
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = input_ready_req_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_val;
  esp_acc_softmax_esp_acc_softmax_mgc_out_dreg_v2 #(.rscid(32'sd5),
  .width(32'sd1)) return_rsci (
      .d(nl_return_rsci_d[0:0]),
      .z(return_rsc_z)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd45),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 #(.rscid(32'sd54)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign input_ready_req_input_ready_req_or_cse = ccs_ccore_start_rsci_idat | (input_ready_req_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_val));
  assign this_rdy_mx0c1 = input_ready_req_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_val & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_rdy <= 1'b0;
    end
    else if ( input_ready_req_input_ready_req_or_cse | this_rdy_mx0c1 ) begin
      this_rdy <= ~ this_rdy_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      input_ready_req_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      input_ready_req_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= input_ready_req_input_ready_req_or_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_bool_Connections_SYN_PORT_Pop
// ------------------------------------------------------------------


module esp_acc_softmax_Connections_Combinational_bool_Connections_SYN_PORT_Pop (
  this_val, this_rdy, this_msg, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  input this_val;
  output this_rdy;
  input this_msg;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_esp_acc_softmax_Connections_Combinational_bool_Connections_SYN_PORT_Pop_core Connections_Combinational_bool_Connections_SYN_PORT_Pop_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> /opt/cad/catapult/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 
  
)( clk,clken,d,q,radr,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" *)
  reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block"
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./softmax_Connections_Combinationalless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_Connections_Combinationalless_boolcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_Connections_Combinationalless_boolcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Sun May  3 17:05:17 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_Connections_Combinational_bool_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_Connections_Combinational_bool_Connections_SYN_PORT_Push_core
    (
  this_val, this_rdy, this_msg, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output this_msg;
  reg this_msg;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg input_ready_ack_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire input_ready_ack_input_ready_ack_or_cse;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = input_ready_ack_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd44),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 #(.rscid(32'sd53)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign input_ready_ack_input_ready_ack_or_cse = ccs_ccore_start_rsci_idat | (input_ready_ack_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_rdy));
  assign this_val_mx0c1 = input_ready_ack_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_val <= 1'b0;
    end
    else if ( input_ready_ack_input_ready_ack_or_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_msg <= 1'b0;
    end
    else if ( (~((~ input_ready_ack_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1)
        | this_rdy)) | ccs_ccore_start_rsci_idat ) begin
      this_msg <= 1'b1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      input_ready_ack_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      input_ready_ack_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= input_ready_ack_input_ready_ack_or_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_bool_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module esp_acc_softmax_Connections_Combinational_bool_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  input this_rdy;
  output this_msg;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_esp_acc_softmax_Connections_Combinational_bool_Connections_SYN_PORT_Push_core Connections_Combinational_bool_Connections_SYN_PORT_Push_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> ./softmax_mgc_shift_l_beh_v5.v 
module esp_acc_softmax_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./softmax_mgc_shift_br_beh_v5.v 
module esp_acc_softmax_mgc_shift_br_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_s(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_s(a,s,1'b0);
     end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshr_u

   //Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction

endmodule

//------> ./softmax_mgc_shift_bl_beh_v5.v 
module esp_acc_softmax_mgc_shift_bl_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate if ( signd_a )
   begin: SGNED
     assign z = fshl_s(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
     assign z = fshl_s(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

endmodule

//------> ./softmax_leading_sign_74_0.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Sun May  3 17:05:19 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_74_0
// ------------------------------------------------------------------


module esp_acc_softmax_leading_sign_74_0 (
  mantissa, rtn
);
  input [73:0] mantissa;
  output [6:0] rtn;


  // Interconnect Declarations
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_24;
  wire c_h_1_27;
  wire c_h_1_28;
  wire c_h_1_29;
  wire c_h_1_30;
  wire c_h_1_33;
  wire c_h_1_34;
  wire c_h_1_35;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc;

  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_1_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_292_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_2_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_or_2_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_nor_nl;

  // Interconnect Declarations for Component Instantiations
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2
      = ~((mantissa[71:70]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1
      = ~((mantissa[73:72]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1
      = ~((mantissa[69:68]!=2'b00));
  assign c_h_1_2 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3
      = (mantissa[67:66]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2
      = ~((mantissa[63:62]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1
      = ~((mantissa[65:64]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1
      = ~((mantissa[61:60]!=2'b00));
  assign c_h_1_5 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4
      = (mantissa[59:58]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1
      & c_h_1_5;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2
      = ~((mantissa[55:54]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1
      = ~((mantissa[57:56]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1
      = ~((mantissa[53:52]!=2'b00));
  assign c_h_1_9 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3
      = (mantissa[51:50]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2
      = ~((mantissa[47:46]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1
      = ~((mantissa[49:48]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1
      = ~((mantissa[45:44]!=2'b00));
  assign c_h_1_12 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5
      = (mantissa[43:42]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1
      & c_h_1_12 & c_h_1_13;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2
      = ~((mantissa[39:38]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1
      = ~((mantissa[41:40]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1
      = ~((mantissa[37:36]!=2'b00));
  assign c_h_1_17 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3
      = (mantissa[35:34]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2
      = ~((mantissa[31:30]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1
      = ~((mantissa[33:32]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1
      = ~((mantissa[29:28]!=2'b00));
  assign c_h_1_20 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4
      = (mantissa[27:26]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1
      & c_h_1_20;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2
      = ~((mantissa[23:22]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1
      = ~((mantissa[25:24]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1
      = ~((mantissa[21:20]!=2'b00));
  assign c_h_1_24 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3
      = (mantissa[19:18]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2
      = ~((mantissa[15:14]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1
      = ~((mantissa[17:16]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1
      = ~((mantissa[13:12]!=2'b00));
  assign c_h_1_27 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2;
  assign c_h_1_28 = c_h_1_24 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3;
  assign c_h_1_29 = c_h_1_21 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_30 = c_h_1_14 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6
      = (mantissa[11:10]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1
      & c_h_1_27 & c_h_1_28 & c_h_1_29;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2
      = ~((mantissa[7:6]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1
      = ~((mantissa[9:8]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1
      = ~((mantissa[5:4]!=2'b00));
  assign c_h_1_33 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3
      = (mantissa[3:2]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1;
  assign c_h_1_34 = c_h_1_33 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3;
  assign c_h_1_35 = c_h_1_30 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc
      = (mantissa[1:0]==2'b00) & c_h_1_34 & c_h_1_35;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_nl
      = c_h_1_30 & (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6);
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_1_nl
      = c_h_1_14 & (c_h_1_29 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5))
      & (~ c_h_1_35);
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_292_nl
      = c_h_1_6 & (c_h_1_13 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4))
      & (~((~(c_h_1_21 & (c_h_1_28 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4))))
      & c_h_1_30)) & (c_h_1_34 | (~ c_h_1_35));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_2_nl
      = c_h_1_2 & (c_h_1_5 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3))
      & (~((~(c_h_1_9 & (c_h_1_12 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~((~(c_h_1_17 & (c_h_1_20 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3))
      & (~((~(c_h_1_24 & (c_h_1_27 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3))))
      & c_h_1_29)))) & c_h_1_30)) & (~((~(c_h_1_33 & (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3)))
      & c_h_1_35));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_or_2_nl
      = (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2))))
      & c_h_1_21)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2))))
      & c_h_1_28)))) & c_h_1_29)))) & c_h_1_30)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2))
      & (~ c_h_1_34))) & c_h_1_35))) | ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_nor_nl
      = ~((mantissa[73]) | (~((mantissa[72:71]!=2'b01))) | (((mantissa[69]) | (~((mantissa[68:67]!=2'b01))))
      & c_h_1_2) | ((~((~((mantissa[65]) | (~((mantissa[64:63]!=2'b01))))) & (~(((mantissa[61])
      | (~((mantissa[60:59]!=2'b01)))) & c_h_1_5)))) & c_h_1_6) | ((~((~((mantissa[57])
      | (~((mantissa[56:55]!=2'b01))))) & (~(((mantissa[53]) | (~((mantissa[52:51]!=2'b01))))
      & c_h_1_9)) & (~((~((~((mantissa[49]) | (~((mantissa[48:47]!=2'b01))))) & (~(((mantissa[45])
      | (~((mantissa[44:43]!=2'b01)))) & c_h_1_12)))) & c_h_1_13)))) & c_h_1_14)
      | ((~((~((mantissa[41]) | (~((mantissa[40:39]!=2'b01))))) & (~(((mantissa[37])
      | (~((mantissa[36:35]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[33]) | (~((mantissa[32:31]!=2'b01)))))
      & (~(((mantissa[29]) | (~((mantissa[28:27]!=2'b01)))) & c_h_1_20)))) & c_h_1_21))
      & (~((~((~((mantissa[25]) | (~((mantissa[24:23]!=2'b01))))) & (~(((mantissa[21])
      | (~((mantissa[20:19]!=2'b01)))) & c_h_1_24)) & (~((~((~((mantissa[17]) | (~((mantissa[16:15]!=2'b01)))))
      & (~(((mantissa[13]) | (~((mantissa[12:11]!=2'b01)))) & c_h_1_27)))) & c_h_1_28))))
      & c_h_1_29)))) & c_h_1_30) | ((~((~((mantissa[9]) | (~((mantissa[8:7]!=2'b01)))))
      & (~(((mantissa[5]) | (~((mantissa[4:3]!=2'b01)))) & c_h_1_33)) & (~((mantissa[1])
      & c_h_1_34)))) & c_h_1_35) | ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc);
  assign rtn = {c_h_1_35 , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_1_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_292_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_2_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_or_2_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_nor_nl};
endmodule




//------> ./softmax_mgc_mul_pipe_beh.v 
//
// File:      $Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v
//
// BASELINE:  Catapult-C version 2006b.63
// MODIFIED:  2007-04-03, tnagler
//
// Note: this file uses Verilog2001 features;
//       please enable Verilog2001 in the flow!

module esp_acc_softmax_mgc_mul_pipe (a, b, clk, en, a_rst, s_rst, z);

    // Parameters:
    parameter integer width_a = 32'd4;  // input a bit width
    parameter         signd_a =  1'b1;  // input a type (1=signed, 0=unsigned)
    parameter integer width_b = 32'd4;  // input b bit width
    parameter         signd_b =  1'b1;  // input b type (1=signed, 0=unsigned)
    parameter integer width_z = 32'd8;  // result bit width (= width_a + width_b)
    parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
    parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
    parameter    a_rst_active =  1'b1;  // unused
    parameter    s_rst_active =  1'b1;  // unused
    parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
    parameter integer n_inreg = 32'd0;  // number of input registers

    localparam integer width_ab = width_a + width_b;  // multiplier result width
    localparam integer n_inreg_min = (n_inreg > 1) ? (n_inreg-1) : 0; // for Synopsys DC

    // I/O ports:
    input  [width_a-1:0] a;      // input A
    input  [width_b-1:0] b;      // input B
    input                clk;    // clock
    input                en;     // enable
    input                a_rst;  // async reset (unused)
    input                s_rst;  // sync reset (unused)
    output [width_z-1:0] z;      // output


    // Input registers:

    wire [width_a-1:0] a_f;
    wire [width_b-1:0] b_f;

    integer i;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(negedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i];
                    b_reg[i+1] <= b_reg[i];
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    else
    begin: POS_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(posedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i];
                    b_reg[i+1] <= b_reg[i];
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    endgenerate


    // Output:
    wire [width_z-1:0]  xz;

    function signed [width_z-1:0] conv_signed;
      input signed [width_ab-1:0] res;
      conv_signed = res[width_z-1:0];
    endfunction

    generate
      wire signed [width_ab-1:0] res;
      if ( (signd_a == 1'b1) && (signd_b == 1'b1) )
      begin: SIGNED_AB
              assign res = $signed(a_f) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b1) && (signd_b == 1'b0) )
      begin: SIGNED_A
              assign res = $signed(a_f) * $signed({1'b0, b_f});
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b0) && (signd_b == 1'b1) )
      begin: SIGNED_B
              assign res = $signed({1'b0,a_f}) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else
      begin: UNSIGNED_AB
              assign res = a_f * b_f;
	      assign xz = res[width_z-1:0];
      end
    endgenerate


    // Output registers:

    reg  [width_z-1:0] reg_array[stages-2:0];
    wire [width_z-1:0] z;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE2
        always @(negedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz;
                else
                    reg_array[i] <= reg_array[i-1];
    end
    else
    begin: POS_EDGE2
        always @(posedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz;
                else
                    reg_array[i] <= reg_array[i-1];
    end
    endgenerate

    assign z = reg_array[stages-2];
endmodule

//------> /opt/cad/catapult/pkgs/ccs_xilinx/hdl/BLOCK_DPRAM_RBW_DUAL.v 
// Memory Type:            BLOCK
// Operating Mode:         True Dual Port (2-Port)
// Clock Mode:             Dual Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_DPRAM_RBW_DUAL
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)

module BLOCK_DPRAM_RBW_DUAL #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 
  
)( adra,adrb,clka,clka_en,clkb,clkb_en,da,db,qa,qb,wea,web);

  input [addr_width-1:0] adra;
  input [addr_width-1:0] adrb;
  input  clka;
  input  clka_en;
  input  clkb;
  input  clkb_en;
  input [data_width-1:0] da;
  input [data_width-1:0] db;
  output [data_width-1:0] qa;
  output [data_width-1:0] qb;
  input  wea;
  input  web;
  
  (* ram_style = "block" *)
  reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block"
  
  reg [data_width-1:0] ramqa;
  reg [data_width-1:0] ramqb;
  
  // Port Map
  // rwA :: ADDRESS adra CLOCK clka ENABLE clka_en DATA_IN da DATA_OUT qa WRITE_ENABLE wea
  // rwB :: ADDRESS adrb CLOCK clkb ENABLE clkb_en DATA_IN db DATA_OUT qb WRITE_ENABLE web

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] adra_reg;
      reg [data_width-1:0] da_reg;
      reg wea_reg;
      reg [addr_width-1:0] adrb_reg;
      reg [data_width-1:0] db_reg;
      reg web_reg;
      
      always @(posedge clka) begin
        if (clka_en) begin
          adra_reg <= adra;
          da_reg <= da;
          wea_reg <= wea;
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
          adrb_reg <= adrb;
          db_reg <= db;
          web_reg <= web;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clka) begin
        if (clka_en) begin
            ramqa <= mem[adra_reg];
            if (wea_reg) begin
              mem[adra_reg] <= da_reg;
            end
        end
      end
      always @(posedge clka) begin
        if (clka_en) begin
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
            ramqb <= mem[adrb_reg];
            if (web_reg) begin
              mem[adrb_reg] <= db_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clka) begin
        if (clka_en) begin
            ramqa <= mem[adra];
            if (wea) begin
              mem[adra] <= da;
            end
        end
      end
      always @(posedge clka) begin
        if (clka_en) begin
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
            ramqb <= mem[adrb];
            if (web) begin
              mem[adrb] <= db;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign qa = ramqa;
      assign qb = ramqb;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpqa;
      reg [data_width-1:0] tmpqb;
      
      always @(posedge clka) begin
        if (clka_en) begin
          tmpqa <= ramqa;
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
          tmpqb <= ramqb;
        end
      end
      
      assign qa = tmpqa;
      assign qb = tmpqb;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1qa;
      reg [data_width-1:0] tmp1qb;
      
      reg [data_width-1:0] tmp2qa;
      reg [data_width-1:0] tmp2qb;
      
      always @(posedge clka) begin
        if (clka_en) begin
          tmp1qa <= ramqa;
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
          tmp1qb <= ramqb;
        end
      end
      
      always @(posedge clka) begin
        if (clka_en) begin
          tmp2qa <= tmp1qa;
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
          tmp2qb <= tmp1qb;
        end
      end
      
      assign qa = tmp2qa;
      assign qb = tmp2qb;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./softmax_Connections_OutBlockingless_sc_dt_sc_bvless_64greater_comma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_Connections_OutBlockingless_sc_dt_sc_bvless_64greater_comma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_Connections_OutBlockingless_sc_dt_sc_bvless_64greater_comma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Sun May  3 17:05:14 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_Connections_OutBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module esp_acc_softmax_esp_acc_softmax_Connections_OutBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Push_core
    (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [63:0] this_msg;
  input [63:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire [63:0] m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [31:0] m_slc_m_31_0_psp_lpi_1_dfm;
  wire and_dcpl;
  reg STORE_OUTPUT_INNER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire STORE_OUTPUT_INNER_LOOP_STORE_OUTPUT_INNER_LOOP_or_cse;
  reg reg_C_32_11011110101011011011111011101111_1_reg_30;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = STORE_OUTPUT_INNER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd7),
  .width(32'sd64)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_in_v1 #(.rscid(32'sd43),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_esp_acc_softmax_ccs_sync_out_vld_v1 #(.rscid(32'sd52)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign this_msg = signext_64_63({reg_C_32_11011110101011011011111011101111_1_reg_30
      , 1'b0 , ({{3{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , reg_C_32_11011110101011011011111011101111_1_reg_30 , 1'b0 , reg_C_32_11011110101011011011111011101111_1_reg_30
      , 1'b0 , ({{1{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{1{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{4{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{2{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{3{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , m_slc_m_31_0_psp_lpi_1_dfm});
  assign STORE_OUTPUT_INNER_LOOP_STORE_OUTPUT_INNER_LOOP_or_cse = ccs_ccore_start_rsci_idat
      | and_dcpl;
  assign and_dcpl = STORE_OUTPUT_INNER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_rdy);
  assign this_val_mx0c1 = STORE_OUTPUT_INNER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_val <= 1'b0;
    end
    else if ( STORE_OUTPUT_INNER_LOOP_STORE_OUTPUT_INNER_LOOP_or_cse | this_val_mx0c1
        ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      reg_C_32_11011110101011011011111011101111_1_reg_30 <= 1'b0;
    end
    else if ( (~((~ STORE_OUTPUT_INNER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1)
        | this_rdy)) | ccs_ccore_start_rsci_idat ) begin
      reg_C_32_11011110101011011011111011101111_1_reg_30 <= 1'b1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      m_slc_m_31_0_psp_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      m_slc_m_31_0_psp_lpi_1_dfm <= m_rsci_idat[31:0];
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      STORE_OUTPUT_INNER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      STORE_OUTPUT_INNER_LOOP_io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= STORE_OUTPUT_INNER_LOOP_STORE_OUTPUT_INNER_LOOP_or_cse;
    end
  end

  function automatic [63:0] signext_64_63;
    input [62:0] vector;
  begin
    signext_64_63= {{1{vector[62]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module esp_acc_softmax_Connections_OutBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  input this_rdy;
  output [63:0] this_msg;
  input [63:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_esp_acc_softmax_Connections_OutBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Push_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_rsc_dat(m_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_ccs_genreg_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_ccs_genreg_v1 (clk, en, arst, srst, d, z);
    parameter integer width   = 1;
    parameter integer ph_clk  = 1;
    parameter integer ph_en   = 1;
    parameter integer ph_arst = 0;
    parameter integer ph_srst = 1;
    parameter         has_en  = 1'b1;

    input clk;
    input en;
    input arst;
    input srst;
    input      [width-1:0] d;
    output reg [width-1:0] z;

    //  Generate parameters
    //  ph_clk | ph_arst | has_en     Label:
    //    1        1          1       GEN_CLK1_ARST1_EN1
    //    1        1          0       GEN_CLK1_ARST1_EN0
    //    1        0          1       GEN_CLK1_ARST0_EN1
    //    1        0          0       GEN_CLK1_ARST0_EN0
    //    0        1          1       GEN_CLK0_ARST1_EN1
    //    0        1          0       GEN_CLK0_ARST1_EN0
    //    0        0          1       GEN_CLK0_ARST0_EN1
    //    0        0          0       GEN_CLK0_ARST0_EN0

    generate
      // Pos edge clock, pos edge async reset, has enable
      if (ph_clk == 1 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK1_ARST1_EN1
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST1_EN1

      // Pos edge clock, pos edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK1_ARST1_EN0
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST1_EN0

      // Pos edge clock, neg edge async reset, has enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK1_ARST0_EN1
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST0_EN1

      // Pos edge clock, neg edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK1_ARST0_EN0
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST0_EN0


      // Neg edge clock, pos edge async reset, has enable
      if (ph_clk == 0 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK0_ARST1_EN1
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST1_EN1

      // Neg edge clock, pos edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK0_ARST1_EN0
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST1_EN0

      // Neg edge clock, neg edge async reset, has enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK0_ARST0_EN1
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST0_EN1

      // Neg edge clock, neg edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK0_ARST0_EN0
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST0_EN0
    endgenerate
endmodule


//------> ./softmax_ccs_fifo_wait_core_v5.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

/*
 *            _________________________________________________
 * WRITER    |                                                 |   READER
 *           |               ccs_fifo_wait_core                |
 *           |             _____________________               |
 *        --<|  din_rdy --<|  ---------------- <|--- dout_rdy <|---
 *           |             |       FIFO         |              |
 *        ---|> din_vld ---|> ----------------  |>-- dout_vld  |>--
 *        ---|>     din ---|> ----------------  |>-- dout      |>--
 *           |             |____________________|              |
 *           |_________________________________________________|
 *
 *    rdy    - can be considered as a notFULL signal
 *    vld    - can be considered as a notEMPTY signal
 *    is_idle - clk can be safely gated
 *
 * Change History:
 *    2019-01-24 - Add assertion to verify rdy signal behavior under reset.
 *                 Fix bug in that behavior.
 */

module esp_acc_softmax_ccs_fifo_wait_core_v5 (clk, en, arst, srst, din_vld, din_rdy, din, dout_vld, dout_rdy, dout, sd, is_idle);

    parameter integer rscid    = 0;     // resource ID
    parameter integer width    = 8;     // fifo width
    parameter integer sz_width = 8;     // size of port for elements in fifo
    parameter integer fifo_sz  = 8;     // fifo depth
    parameter integer ph_clk   = 1;  // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1;  // clock enable polarity
    parameter integer ph_arst  = 1;  // async reset polarity
    parameter integer ph_srst  = 1;  // sync reset polarity
    parameter integer ph_log2  = 3;     // log2(fifo_sz)

    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 din_vld;    // writer has valid data
    output                din_rdy;    // fifo ready for data (not full)
    input  [width-1:0]    din;
    output                dout_vld;   // fifo has valid data (not empty)
    input                 dout_rdy;   // reader ready for data
    output [width-1:0]    dout;
    output [sz_width-1:0] sd;
    output                is_idle;

    localparam integer fifo_b  = width * fifo_sz;
    localparam integer fifo_mx = (fifo_sz > 0) ? (fifo_sz-1) : 0 ;
    localparam integer fifo_mx_over_8 = fifo_mx / 8 ;

    reg      [fifo_mx:0] stat_pre;
    wire     [fifo_mx:0] stat;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    wire     [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    reg      [fifo_mx:0] en_l;
    reg      [fifo_mx_over_8:0] en_l_s;

    reg      [width-1:0] buff_nxt;

    reg                  stat_nxt;
    reg                  stat_behind;
    reg                  stat_ahead;
    reg                  en_l_var;

    integer              i;
    genvar               eni;

    wire [32:0]          size_t;
    reg  [31:0]          count;
    reg  [31:0]          count_t;
    reg  [32:0]          n_elem;
// synopsys translate_off
    reg  [31:0]          peak;
    initial
    begin
      count = 32'b0;
      peak  = 32'b0;
    end
// synopsys translate_on
  wire din_rdy_drv  ;
  wire dout_vld_drv ;
    wire                 active;
    wire                 din_vld_int;
    wire                 hs_init;

    //assign din_rdy  = din_rdy_drv;    // dout_rdy | (~stat[0] & hs_init);   // original
    assign din_rdy = (fifo_sz > 0) ? (~stat[0] | dout_rdy) && hs_init : dout_rdy ;
    assign dout_vld = dout_vld_drv;
    assign is_idle = (~((din_vld && din_rdy) || (dout_vld && dout_rdy))) && hs_init;

    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
    assign din_vld_int = din_vld & hs_init;
    assign active =   (din_vld_int & din_rdy_drv) | (dout_rdy & dout_vld_drv);

      assign din_rdy_drv = dout_rdy | (~stat[0] & hs_init);
      assign dout_vld_drv = din_vld_int | stat[fifo_sz-1];

      assign size_t = (count - {31'b0 , (dout_rdy & stat[fifo_sz-1])}) + { 31'b0, din_vld_int};
      assign sd = size_t[sz_width-1:0];

      assign dout = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : din;

      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          stat_behind = (i != 0) ? stat[i-1] : 1'b0;
          stat_ahead  = (i != (fifo_sz-1)) ? stat[i+1] : 1'b1;

          // Determine if this buffer element will have data
          stat_nxt = stat_ahead &                       // valid element ahead of this one (or head)
                       (stat_behind                     // valid element behind this one
                         | (stat[i] & (~dout_rdy))      // valid element and output not ready (in use, no tx)
                         | (stat[i] & din_vld_int)      // valid element and input has data
                         | (din_vld_int  & (~dout_rdy)) // input has data and output not ready
                       );
          stat_pre[i] = stat_nxt;

          if (dout_rdy & stat_behind )
          begin
            // pop n shift
            buff_nxt[0+:width] = buff[width*(i-1)+:width];
            en_l_var = 1'b1;
          end
          else if (din_vld_int & stat_nxt & ~((~dout_rdy) & stat[i]))
          begin
            // update tail with input data
            buff_nxt = din;
            en_l_var = 1'b1;
          end
          else
          begin
            // no-op, disable register
            buff_nxt = din; // Don't care input to disabled flop
            en_l_var = 1'b0;
          end
          buff_pre[width*i+:width] = buff_nxt[0+:width];

          if (ph_en != 0)
            en_l[i] = en & en_l_var;
          else
            en_l[i] = en | ~en_l_var;

          if ((stat_ahead == 1'b1) & (stat[i] == 1'b0))
            //found tail, update the number of elements for count
            n_elem = ($unsigned(fifo_sz) - 1) - $unsigned(i);
        end //for loop

        // Enable for stat registers (partitioned into banks of eight)
        // Take care of the head first
        if (ph_en != 0)
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en & active;
        else
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en | ~active;

        // Now every eight
        for (i = fifo_sz-1; i >= 7; i = i - 1)
        begin
          if (($unsigned(i)%8) == 0)
          begin
            if (ph_en != 0)
              en_l_s[(i/8)-1] = en & (stat[i]) & (active);
            else
              en_l_s[(i/8)-1] = en | ~(stat[i]) | ~(active);
          end
        end

        // Update count and peak
        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = fifo_sz;
        else
          count_t = n_elem[31:0];
        count = count_t;
// synopsys translate_off
        if ( peak < count )
          peak = count;
// synopsys translate_on
      end //FIFOPROC

      // Handshake valid after reset
      esp_acc_softmax_ccs_genreg_v1
      #(
        .width   (1),
        .ph_clk  (ph_clk),
        .ph_en   (1),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .has_en  (1'b0)
      )
      HS_INIT_REG
      (
        .clk     (clk),
        .en      (1'b1),
        .arst    (arst),
        .srst    (srst),
        .d       (1'b1),
        .z       (hs_init)
      );

      // Buffer and status registers
      for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
      begin: GEN_REGS
        esp_acc_softmax_ccs_genreg_v1
        #(
          .width   (1),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        STATREG
        (
          .clk     (clk),
          .en      (en_l_s[eni/8]),
          .arst    (arst),
          .srst    (srst),
          .d       (stat_pre[eni]),
          .z       (stat[eni])
        );

        esp_acc_softmax_ccs_genreg_v1
        #(
          .width   (width),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        BUFREG
        (
          .clk     (clk),
          .en      (en_l[eni]),
          .arst    (arst),
          .srst    (srst),
          .d       (buff_pre[width*eni+:width]),
          .z       (buff[width*eni+:width])
        );
      end

    end
    else
    begin: FEED_THRU
      assign din_rdy_drv  = dout_rdy;
      assign dout_vld_drv = din_vld;
      assign dout     = din;
      // non-blocking is not II=1 when fifo_sz=0
      assign sd = {{(sz_width-1){1'b0}}, (din_vld & ~dout_rdy)};
    end
    endgenerate

`ifdef RDY_ASRT
    generate
    if (ph_clk==1)
    begin: POS_CLK_ASSERT

       property rdyAsrt ;
         @(posedge clk) ((srst==ph_srst) || (arst==ph_arst)) |=> (din_rdy==0);
       endproperty
       a1Pos: assert property(rdyAsrt);

    end else if (ph_clk==0)
    begin: NEG_CLK_ASSERT

       property rdyAsrt ;
         @(negedge clk) ((srst==ph_srst) || (arst==ph_arst)) |=> (din_rdy==0);
       endproperty
       a1Neg: assert property(rdyAsrt);

    end
    endgenerate

`endif

endmodule



//------> ./softmax_ccs_pipe_v5.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
/*
 *
 *            _______________________________________________
 * WRITER    |                                              |          READER
 *           |                 ccs_pipe                     |
 *           |            ______________________            |
 *        --<| din_rdy --<|  ---------------- <|---dout_rdy<|---
 *           |            |       FIFO         |            |
 *        ---|>din_vld ---|> ----------------  |>--dout_vld |>--
 *        ---|>din -------|> ----------------  |> -----dout |>--
 *           |            |____________________|            |
 *           |______________________________________________|
 *
 *    din_rdy     - can be considered as a notFULL signal
 *    dout_vld    - can be considered as a notEMPTY signal
 *    write_stall - an internal debug signal formed from din_vld & !din_rdy
 *    read_stall  - an internal debug signal formed from dout_rdy & !dout_vld
 *    is_idle     - indicates the clock can be safely gated
 */

module esp_acc_softmax_ccs_pipe_v5 (clk, en, arst, srst, din_rdy, din_vld, din, dout_rdy, dout_vld, dout, sz, sz_req, is_idle);

    parameter integer rscid    = 0; // resource ID
    parameter integer width    = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz  = 8; // fifo depth
    parameter integer log2_sz  = 3; // log2(fifo_sz)
    parameter integer ph_clk   = 1; // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1; // clock enable polarity
    parameter integer ph_arst  = 1; // async reset polarity
    parameter integer ph_srst  = 1; // sync reset polarity

    // clock
    input              clk;
    input              en;
    input              arst;
    input              srst;

    // writer
    output             din_rdy;
    input              din_vld;
    input  [width-1:0] din;

    // reader
    input              dout_rdy;
    output             dout_vld;
    output [width-1:0] dout;

    // size
    output [sz_width-1:0] sz;
    input                 sz_req;
    output                is_idle;

// synopsys translate_off
    wire   write_stall;
    wire   read_stall;
    assign write_stall = din_vld & !din_rdy;
    assign read_stall  = dout_rdy & !dout_vld;
// synopsys translate_on

    esp_acc_softmax_ccs_fifo_wait_core_v5
    #(
        .rscid    (rscid),
        .width    (width),
        .sz_width (sz_width),
        .fifo_sz  (fifo_sz),
        .ph_clk   (ph_clk),
        .ph_en    (ph_en),
        .ph_arst  (ph_arst),
        .ph_srst  (ph_srst),
        .ph_log2  (log2_sz)
    )
    FIFO
    (
        .clk      (clk),
        .en       (en),
        .arst     (arst),
        .srst     (srst),
        .din_vld  (din_vld),
        .din_rdy  (din_rdy),
        .din      (din),
        .dout_vld (dout_vld),
        .dout_rdy (dout_rdy),
        .dout     (dout),
        .sd       (sz),
        .is_idle  (is_idle)
    );

endmodule


//------> ./softmax.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Sun May  3 17:06:21 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_20_7_32_128_128_32_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_20_7_32_128_128_32_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [31:0] q;
  output [6:0] radr;
  output we;
  output [31:0] d;
  output [6:0] wadr;
  input clken_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_store_output_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_store_output_fsm (
  clk, rst, store_output_wen, fsm_output, WAIT_FOR_CONFIG_LOOP_C_0_tr0, store_output_rlp_C_0_tr0,
      COMPUTE_BATCH_LOOP_C_0_tr0, STORE_OUTPUT_INNER_LOOP_C_0_tr0, STORE_MAIN_LOOP_C_130_tr0,
      COMPUTE_BATCH_LOOP_C_1_tr0
);
  input clk;
  input rst;
  input store_output_wen;
  output [7:0] fsm_output;
  reg [7:0] fsm_output;
  input WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  input store_output_rlp_C_0_tr0;
  input COMPUTE_BATCH_LOOP_C_0_tr0;
  input STORE_OUTPUT_INNER_LOOP_C_0_tr0;
  input STORE_MAIN_LOOP_C_130_tr0;
  input COMPUTE_BATCH_LOOP_C_1_tr0;


  // FSM State Type Declaration for esp_acc_softmax_softmax_store_output_store_output_store_output_fsm_1
  parameter
    WAIT_FOR_CONFIG_LOOP_C_0 = 8'd0,
    store_output_rlp_C_0 = 8'd1,
    COMPUTE_BATCH_LOOP_C_0 = 8'd2,
    STORE_MAIN_LOOP_C_0 = 8'd3,
    STORE_MAIN_LOOP_C_1 = 8'd4,
    STORE_MAIN_LOOP_C_2 = 8'd5,
    STORE_MAIN_LOOP_C_3 = 8'd6,
    STORE_MAIN_LOOP_C_4 = 8'd7,
    STORE_MAIN_LOOP_C_5 = 8'd8,
    STORE_MAIN_LOOP_C_6 = 8'd9,
    STORE_MAIN_LOOP_C_7 = 8'd10,
    STORE_MAIN_LOOP_C_8 = 8'd11,
    STORE_MAIN_LOOP_C_9 = 8'd12,
    STORE_MAIN_LOOP_C_10 = 8'd13,
    STORE_MAIN_LOOP_C_11 = 8'd14,
    STORE_MAIN_LOOP_C_12 = 8'd15,
    STORE_MAIN_LOOP_C_13 = 8'd16,
    STORE_MAIN_LOOP_C_14 = 8'd17,
    STORE_MAIN_LOOP_C_15 = 8'd18,
    STORE_MAIN_LOOP_C_16 = 8'd19,
    STORE_MAIN_LOOP_C_17 = 8'd20,
    STORE_MAIN_LOOP_C_18 = 8'd21,
    STORE_MAIN_LOOP_C_19 = 8'd22,
    STORE_MAIN_LOOP_C_20 = 8'd23,
    STORE_MAIN_LOOP_C_21 = 8'd24,
    STORE_MAIN_LOOP_C_22 = 8'd25,
    STORE_MAIN_LOOP_C_23 = 8'd26,
    STORE_MAIN_LOOP_C_24 = 8'd27,
    STORE_MAIN_LOOP_C_25 = 8'd28,
    STORE_MAIN_LOOP_C_26 = 8'd29,
    STORE_MAIN_LOOP_C_27 = 8'd30,
    STORE_MAIN_LOOP_C_28 = 8'd31,
    STORE_MAIN_LOOP_C_29 = 8'd32,
    STORE_MAIN_LOOP_C_30 = 8'd33,
    STORE_MAIN_LOOP_C_31 = 8'd34,
    STORE_MAIN_LOOP_C_32 = 8'd35,
    STORE_MAIN_LOOP_C_33 = 8'd36,
    STORE_MAIN_LOOP_C_34 = 8'd37,
    STORE_MAIN_LOOP_C_35 = 8'd38,
    STORE_MAIN_LOOP_C_36 = 8'd39,
    STORE_MAIN_LOOP_C_37 = 8'd40,
    STORE_MAIN_LOOP_C_38 = 8'd41,
    STORE_MAIN_LOOP_C_39 = 8'd42,
    STORE_MAIN_LOOP_C_40 = 8'd43,
    STORE_MAIN_LOOP_C_41 = 8'd44,
    STORE_MAIN_LOOP_C_42 = 8'd45,
    STORE_MAIN_LOOP_C_43 = 8'd46,
    STORE_MAIN_LOOP_C_44 = 8'd47,
    STORE_MAIN_LOOP_C_45 = 8'd48,
    STORE_MAIN_LOOP_C_46 = 8'd49,
    STORE_MAIN_LOOP_C_47 = 8'd50,
    STORE_MAIN_LOOP_C_48 = 8'd51,
    STORE_MAIN_LOOP_C_49 = 8'd52,
    STORE_MAIN_LOOP_C_50 = 8'd53,
    STORE_MAIN_LOOP_C_51 = 8'd54,
    STORE_MAIN_LOOP_C_52 = 8'd55,
    STORE_MAIN_LOOP_C_53 = 8'd56,
    STORE_MAIN_LOOP_C_54 = 8'd57,
    STORE_MAIN_LOOP_C_55 = 8'd58,
    STORE_MAIN_LOOP_C_56 = 8'd59,
    STORE_MAIN_LOOP_C_57 = 8'd60,
    STORE_MAIN_LOOP_C_58 = 8'd61,
    STORE_MAIN_LOOP_C_59 = 8'd62,
    STORE_MAIN_LOOP_C_60 = 8'd63,
    STORE_MAIN_LOOP_C_61 = 8'd64,
    STORE_MAIN_LOOP_C_62 = 8'd65,
    STORE_MAIN_LOOP_C_63 = 8'd66,
    STORE_MAIN_LOOP_C_64 = 8'd67,
    STORE_MAIN_LOOP_C_65 = 8'd68,
    STORE_MAIN_LOOP_C_66 = 8'd69,
    STORE_MAIN_LOOP_C_67 = 8'd70,
    STORE_MAIN_LOOP_C_68 = 8'd71,
    STORE_MAIN_LOOP_C_69 = 8'd72,
    STORE_MAIN_LOOP_C_70 = 8'd73,
    STORE_MAIN_LOOP_C_71 = 8'd74,
    STORE_MAIN_LOOP_C_72 = 8'd75,
    STORE_MAIN_LOOP_C_73 = 8'd76,
    STORE_MAIN_LOOP_C_74 = 8'd77,
    STORE_MAIN_LOOP_C_75 = 8'd78,
    STORE_MAIN_LOOP_C_76 = 8'd79,
    STORE_MAIN_LOOP_C_77 = 8'd80,
    STORE_MAIN_LOOP_C_78 = 8'd81,
    STORE_MAIN_LOOP_C_79 = 8'd82,
    STORE_MAIN_LOOP_C_80 = 8'd83,
    STORE_MAIN_LOOP_C_81 = 8'd84,
    STORE_MAIN_LOOP_C_82 = 8'd85,
    STORE_MAIN_LOOP_C_83 = 8'd86,
    STORE_MAIN_LOOP_C_84 = 8'd87,
    STORE_MAIN_LOOP_C_85 = 8'd88,
    STORE_MAIN_LOOP_C_86 = 8'd89,
    STORE_MAIN_LOOP_C_87 = 8'd90,
    STORE_MAIN_LOOP_C_88 = 8'd91,
    STORE_MAIN_LOOP_C_89 = 8'd92,
    STORE_MAIN_LOOP_C_90 = 8'd93,
    STORE_MAIN_LOOP_C_91 = 8'd94,
    STORE_MAIN_LOOP_C_92 = 8'd95,
    STORE_MAIN_LOOP_C_93 = 8'd96,
    STORE_MAIN_LOOP_C_94 = 8'd97,
    STORE_MAIN_LOOP_C_95 = 8'd98,
    STORE_MAIN_LOOP_C_96 = 8'd99,
    STORE_MAIN_LOOP_C_97 = 8'd100,
    STORE_MAIN_LOOP_C_98 = 8'd101,
    STORE_MAIN_LOOP_C_99 = 8'd102,
    STORE_MAIN_LOOP_C_100 = 8'd103,
    STORE_MAIN_LOOP_C_101 = 8'd104,
    STORE_MAIN_LOOP_C_102 = 8'd105,
    STORE_MAIN_LOOP_C_103 = 8'd106,
    STORE_MAIN_LOOP_C_104 = 8'd107,
    STORE_MAIN_LOOP_C_105 = 8'd108,
    STORE_MAIN_LOOP_C_106 = 8'd109,
    STORE_MAIN_LOOP_C_107 = 8'd110,
    STORE_MAIN_LOOP_C_108 = 8'd111,
    STORE_MAIN_LOOP_C_109 = 8'd112,
    STORE_MAIN_LOOP_C_110 = 8'd113,
    STORE_MAIN_LOOP_C_111 = 8'd114,
    STORE_MAIN_LOOP_C_112 = 8'd115,
    STORE_MAIN_LOOP_C_113 = 8'd116,
    STORE_MAIN_LOOP_C_114 = 8'd117,
    STORE_MAIN_LOOP_C_115 = 8'd118,
    STORE_MAIN_LOOP_C_116 = 8'd119,
    STORE_MAIN_LOOP_C_117 = 8'd120,
    STORE_MAIN_LOOP_C_118 = 8'd121,
    STORE_MAIN_LOOP_C_119 = 8'd122,
    STORE_MAIN_LOOP_C_120 = 8'd123,
    STORE_MAIN_LOOP_C_121 = 8'd124,
    STORE_MAIN_LOOP_C_122 = 8'd125,
    STORE_MAIN_LOOP_C_123 = 8'd126,
    STORE_MAIN_LOOP_C_124 = 8'd127,
    STORE_MAIN_LOOP_C_125 = 8'd128,
    STORE_MAIN_LOOP_C_126 = 8'd129,
    STORE_MAIN_LOOP_C_127 = 8'd130,
    STORE_MAIN_LOOP_C_128 = 8'd131,
    STORE_MAIN_LOOP_C_129 = 8'd132,
    STORE_OUTPUT_INNER_LOOP_C_0 = 8'd133,
    STORE_MAIN_LOOP_C_130 = 8'd134,
    COMPUTE_BATCH_LOOP_C_1 = 8'd135,
    store_output_rlp_C_1 = 8'd136,
    PROCESS_DONE_LOOP_C_0 = 8'd137;

  reg [7:0] state_var;
  reg [7:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_softmax_softmax_store_output_store_output_store_output_fsm_1
    case (state_var)
      store_output_rlp_C_0 : begin
        fsm_output = 8'b00000001;
        if ( store_output_rlp_C_0_tr0 ) begin
          state_var_NS = COMPUTE_BATCH_LOOP_C_0;
        end
        else begin
          state_var_NS = store_output_rlp_C_1;
        end
      end
      COMPUTE_BATCH_LOOP_C_0 : begin
        fsm_output = 8'b00000010;
        if ( COMPUTE_BATCH_LOOP_C_0_tr0 ) begin
          state_var_NS = COMPUTE_BATCH_LOOP_C_1;
        end
        else begin
          state_var_NS = STORE_MAIN_LOOP_C_0;
        end
      end
      STORE_MAIN_LOOP_C_0 : begin
        fsm_output = 8'b00000011;
        state_var_NS = STORE_MAIN_LOOP_C_1;
      end
      STORE_MAIN_LOOP_C_1 : begin
        fsm_output = 8'b00000100;
        state_var_NS = STORE_MAIN_LOOP_C_2;
      end
      STORE_MAIN_LOOP_C_2 : begin
        fsm_output = 8'b00000101;
        state_var_NS = STORE_MAIN_LOOP_C_3;
      end
      STORE_MAIN_LOOP_C_3 : begin
        fsm_output = 8'b00000110;
        state_var_NS = STORE_MAIN_LOOP_C_4;
      end
      STORE_MAIN_LOOP_C_4 : begin
        fsm_output = 8'b00000111;
        state_var_NS = STORE_MAIN_LOOP_C_5;
      end
      STORE_MAIN_LOOP_C_5 : begin
        fsm_output = 8'b00001000;
        state_var_NS = STORE_MAIN_LOOP_C_6;
      end
      STORE_MAIN_LOOP_C_6 : begin
        fsm_output = 8'b00001001;
        state_var_NS = STORE_MAIN_LOOP_C_7;
      end
      STORE_MAIN_LOOP_C_7 : begin
        fsm_output = 8'b00001010;
        state_var_NS = STORE_MAIN_LOOP_C_8;
      end
      STORE_MAIN_LOOP_C_8 : begin
        fsm_output = 8'b00001011;
        state_var_NS = STORE_MAIN_LOOP_C_9;
      end
      STORE_MAIN_LOOP_C_9 : begin
        fsm_output = 8'b00001100;
        state_var_NS = STORE_MAIN_LOOP_C_10;
      end
      STORE_MAIN_LOOP_C_10 : begin
        fsm_output = 8'b00001101;
        state_var_NS = STORE_MAIN_LOOP_C_11;
      end
      STORE_MAIN_LOOP_C_11 : begin
        fsm_output = 8'b00001110;
        state_var_NS = STORE_MAIN_LOOP_C_12;
      end
      STORE_MAIN_LOOP_C_12 : begin
        fsm_output = 8'b00001111;
        state_var_NS = STORE_MAIN_LOOP_C_13;
      end
      STORE_MAIN_LOOP_C_13 : begin
        fsm_output = 8'b00010000;
        state_var_NS = STORE_MAIN_LOOP_C_14;
      end
      STORE_MAIN_LOOP_C_14 : begin
        fsm_output = 8'b00010001;
        state_var_NS = STORE_MAIN_LOOP_C_15;
      end
      STORE_MAIN_LOOP_C_15 : begin
        fsm_output = 8'b00010010;
        state_var_NS = STORE_MAIN_LOOP_C_16;
      end
      STORE_MAIN_LOOP_C_16 : begin
        fsm_output = 8'b00010011;
        state_var_NS = STORE_MAIN_LOOP_C_17;
      end
      STORE_MAIN_LOOP_C_17 : begin
        fsm_output = 8'b00010100;
        state_var_NS = STORE_MAIN_LOOP_C_18;
      end
      STORE_MAIN_LOOP_C_18 : begin
        fsm_output = 8'b00010101;
        state_var_NS = STORE_MAIN_LOOP_C_19;
      end
      STORE_MAIN_LOOP_C_19 : begin
        fsm_output = 8'b00010110;
        state_var_NS = STORE_MAIN_LOOP_C_20;
      end
      STORE_MAIN_LOOP_C_20 : begin
        fsm_output = 8'b00010111;
        state_var_NS = STORE_MAIN_LOOP_C_21;
      end
      STORE_MAIN_LOOP_C_21 : begin
        fsm_output = 8'b00011000;
        state_var_NS = STORE_MAIN_LOOP_C_22;
      end
      STORE_MAIN_LOOP_C_22 : begin
        fsm_output = 8'b00011001;
        state_var_NS = STORE_MAIN_LOOP_C_23;
      end
      STORE_MAIN_LOOP_C_23 : begin
        fsm_output = 8'b00011010;
        state_var_NS = STORE_MAIN_LOOP_C_24;
      end
      STORE_MAIN_LOOP_C_24 : begin
        fsm_output = 8'b00011011;
        state_var_NS = STORE_MAIN_LOOP_C_25;
      end
      STORE_MAIN_LOOP_C_25 : begin
        fsm_output = 8'b00011100;
        state_var_NS = STORE_MAIN_LOOP_C_26;
      end
      STORE_MAIN_LOOP_C_26 : begin
        fsm_output = 8'b00011101;
        state_var_NS = STORE_MAIN_LOOP_C_27;
      end
      STORE_MAIN_LOOP_C_27 : begin
        fsm_output = 8'b00011110;
        state_var_NS = STORE_MAIN_LOOP_C_28;
      end
      STORE_MAIN_LOOP_C_28 : begin
        fsm_output = 8'b00011111;
        state_var_NS = STORE_MAIN_LOOP_C_29;
      end
      STORE_MAIN_LOOP_C_29 : begin
        fsm_output = 8'b00100000;
        state_var_NS = STORE_MAIN_LOOP_C_30;
      end
      STORE_MAIN_LOOP_C_30 : begin
        fsm_output = 8'b00100001;
        state_var_NS = STORE_MAIN_LOOP_C_31;
      end
      STORE_MAIN_LOOP_C_31 : begin
        fsm_output = 8'b00100010;
        state_var_NS = STORE_MAIN_LOOP_C_32;
      end
      STORE_MAIN_LOOP_C_32 : begin
        fsm_output = 8'b00100011;
        state_var_NS = STORE_MAIN_LOOP_C_33;
      end
      STORE_MAIN_LOOP_C_33 : begin
        fsm_output = 8'b00100100;
        state_var_NS = STORE_MAIN_LOOP_C_34;
      end
      STORE_MAIN_LOOP_C_34 : begin
        fsm_output = 8'b00100101;
        state_var_NS = STORE_MAIN_LOOP_C_35;
      end
      STORE_MAIN_LOOP_C_35 : begin
        fsm_output = 8'b00100110;
        state_var_NS = STORE_MAIN_LOOP_C_36;
      end
      STORE_MAIN_LOOP_C_36 : begin
        fsm_output = 8'b00100111;
        state_var_NS = STORE_MAIN_LOOP_C_37;
      end
      STORE_MAIN_LOOP_C_37 : begin
        fsm_output = 8'b00101000;
        state_var_NS = STORE_MAIN_LOOP_C_38;
      end
      STORE_MAIN_LOOP_C_38 : begin
        fsm_output = 8'b00101001;
        state_var_NS = STORE_MAIN_LOOP_C_39;
      end
      STORE_MAIN_LOOP_C_39 : begin
        fsm_output = 8'b00101010;
        state_var_NS = STORE_MAIN_LOOP_C_40;
      end
      STORE_MAIN_LOOP_C_40 : begin
        fsm_output = 8'b00101011;
        state_var_NS = STORE_MAIN_LOOP_C_41;
      end
      STORE_MAIN_LOOP_C_41 : begin
        fsm_output = 8'b00101100;
        state_var_NS = STORE_MAIN_LOOP_C_42;
      end
      STORE_MAIN_LOOP_C_42 : begin
        fsm_output = 8'b00101101;
        state_var_NS = STORE_MAIN_LOOP_C_43;
      end
      STORE_MAIN_LOOP_C_43 : begin
        fsm_output = 8'b00101110;
        state_var_NS = STORE_MAIN_LOOP_C_44;
      end
      STORE_MAIN_LOOP_C_44 : begin
        fsm_output = 8'b00101111;
        state_var_NS = STORE_MAIN_LOOP_C_45;
      end
      STORE_MAIN_LOOP_C_45 : begin
        fsm_output = 8'b00110000;
        state_var_NS = STORE_MAIN_LOOP_C_46;
      end
      STORE_MAIN_LOOP_C_46 : begin
        fsm_output = 8'b00110001;
        state_var_NS = STORE_MAIN_LOOP_C_47;
      end
      STORE_MAIN_LOOP_C_47 : begin
        fsm_output = 8'b00110010;
        state_var_NS = STORE_MAIN_LOOP_C_48;
      end
      STORE_MAIN_LOOP_C_48 : begin
        fsm_output = 8'b00110011;
        state_var_NS = STORE_MAIN_LOOP_C_49;
      end
      STORE_MAIN_LOOP_C_49 : begin
        fsm_output = 8'b00110100;
        state_var_NS = STORE_MAIN_LOOP_C_50;
      end
      STORE_MAIN_LOOP_C_50 : begin
        fsm_output = 8'b00110101;
        state_var_NS = STORE_MAIN_LOOP_C_51;
      end
      STORE_MAIN_LOOP_C_51 : begin
        fsm_output = 8'b00110110;
        state_var_NS = STORE_MAIN_LOOP_C_52;
      end
      STORE_MAIN_LOOP_C_52 : begin
        fsm_output = 8'b00110111;
        state_var_NS = STORE_MAIN_LOOP_C_53;
      end
      STORE_MAIN_LOOP_C_53 : begin
        fsm_output = 8'b00111000;
        state_var_NS = STORE_MAIN_LOOP_C_54;
      end
      STORE_MAIN_LOOP_C_54 : begin
        fsm_output = 8'b00111001;
        state_var_NS = STORE_MAIN_LOOP_C_55;
      end
      STORE_MAIN_LOOP_C_55 : begin
        fsm_output = 8'b00111010;
        state_var_NS = STORE_MAIN_LOOP_C_56;
      end
      STORE_MAIN_LOOP_C_56 : begin
        fsm_output = 8'b00111011;
        state_var_NS = STORE_MAIN_LOOP_C_57;
      end
      STORE_MAIN_LOOP_C_57 : begin
        fsm_output = 8'b00111100;
        state_var_NS = STORE_MAIN_LOOP_C_58;
      end
      STORE_MAIN_LOOP_C_58 : begin
        fsm_output = 8'b00111101;
        state_var_NS = STORE_MAIN_LOOP_C_59;
      end
      STORE_MAIN_LOOP_C_59 : begin
        fsm_output = 8'b00111110;
        state_var_NS = STORE_MAIN_LOOP_C_60;
      end
      STORE_MAIN_LOOP_C_60 : begin
        fsm_output = 8'b00111111;
        state_var_NS = STORE_MAIN_LOOP_C_61;
      end
      STORE_MAIN_LOOP_C_61 : begin
        fsm_output = 8'b01000000;
        state_var_NS = STORE_MAIN_LOOP_C_62;
      end
      STORE_MAIN_LOOP_C_62 : begin
        fsm_output = 8'b01000001;
        state_var_NS = STORE_MAIN_LOOP_C_63;
      end
      STORE_MAIN_LOOP_C_63 : begin
        fsm_output = 8'b01000010;
        state_var_NS = STORE_MAIN_LOOP_C_64;
      end
      STORE_MAIN_LOOP_C_64 : begin
        fsm_output = 8'b01000011;
        state_var_NS = STORE_MAIN_LOOP_C_65;
      end
      STORE_MAIN_LOOP_C_65 : begin
        fsm_output = 8'b01000100;
        state_var_NS = STORE_MAIN_LOOP_C_66;
      end
      STORE_MAIN_LOOP_C_66 : begin
        fsm_output = 8'b01000101;
        state_var_NS = STORE_MAIN_LOOP_C_67;
      end
      STORE_MAIN_LOOP_C_67 : begin
        fsm_output = 8'b01000110;
        state_var_NS = STORE_MAIN_LOOP_C_68;
      end
      STORE_MAIN_LOOP_C_68 : begin
        fsm_output = 8'b01000111;
        state_var_NS = STORE_MAIN_LOOP_C_69;
      end
      STORE_MAIN_LOOP_C_69 : begin
        fsm_output = 8'b01001000;
        state_var_NS = STORE_MAIN_LOOP_C_70;
      end
      STORE_MAIN_LOOP_C_70 : begin
        fsm_output = 8'b01001001;
        state_var_NS = STORE_MAIN_LOOP_C_71;
      end
      STORE_MAIN_LOOP_C_71 : begin
        fsm_output = 8'b01001010;
        state_var_NS = STORE_MAIN_LOOP_C_72;
      end
      STORE_MAIN_LOOP_C_72 : begin
        fsm_output = 8'b01001011;
        state_var_NS = STORE_MAIN_LOOP_C_73;
      end
      STORE_MAIN_LOOP_C_73 : begin
        fsm_output = 8'b01001100;
        state_var_NS = STORE_MAIN_LOOP_C_74;
      end
      STORE_MAIN_LOOP_C_74 : begin
        fsm_output = 8'b01001101;
        state_var_NS = STORE_MAIN_LOOP_C_75;
      end
      STORE_MAIN_LOOP_C_75 : begin
        fsm_output = 8'b01001110;
        state_var_NS = STORE_MAIN_LOOP_C_76;
      end
      STORE_MAIN_LOOP_C_76 : begin
        fsm_output = 8'b01001111;
        state_var_NS = STORE_MAIN_LOOP_C_77;
      end
      STORE_MAIN_LOOP_C_77 : begin
        fsm_output = 8'b01010000;
        state_var_NS = STORE_MAIN_LOOP_C_78;
      end
      STORE_MAIN_LOOP_C_78 : begin
        fsm_output = 8'b01010001;
        state_var_NS = STORE_MAIN_LOOP_C_79;
      end
      STORE_MAIN_LOOP_C_79 : begin
        fsm_output = 8'b01010010;
        state_var_NS = STORE_MAIN_LOOP_C_80;
      end
      STORE_MAIN_LOOP_C_80 : begin
        fsm_output = 8'b01010011;
        state_var_NS = STORE_MAIN_LOOP_C_81;
      end
      STORE_MAIN_LOOP_C_81 : begin
        fsm_output = 8'b01010100;
        state_var_NS = STORE_MAIN_LOOP_C_82;
      end
      STORE_MAIN_LOOP_C_82 : begin
        fsm_output = 8'b01010101;
        state_var_NS = STORE_MAIN_LOOP_C_83;
      end
      STORE_MAIN_LOOP_C_83 : begin
        fsm_output = 8'b01010110;
        state_var_NS = STORE_MAIN_LOOP_C_84;
      end
      STORE_MAIN_LOOP_C_84 : begin
        fsm_output = 8'b01010111;
        state_var_NS = STORE_MAIN_LOOP_C_85;
      end
      STORE_MAIN_LOOP_C_85 : begin
        fsm_output = 8'b01011000;
        state_var_NS = STORE_MAIN_LOOP_C_86;
      end
      STORE_MAIN_LOOP_C_86 : begin
        fsm_output = 8'b01011001;
        state_var_NS = STORE_MAIN_LOOP_C_87;
      end
      STORE_MAIN_LOOP_C_87 : begin
        fsm_output = 8'b01011010;
        state_var_NS = STORE_MAIN_LOOP_C_88;
      end
      STORE_MAIN_LOOP_C_88 : begin
        fsm_output = 8'b01011011;
        state_var_NS = STORE_MAIN_LOOP_C_89;
      end
      STORE_MAIN_LOOP_C_89 : begin
        fsm_output = 8'b01011100;
        state_var_NS = STORE_MAIN_LOOP_C_90;
      end
      STORE_MAIN_LOOP_C_90 : begin
        fsm_output = 8'b01011101;
        state_var_NS = STORE_MAIN_LOOP_C_91;
      end
      STORE_MAIN_LOOP_C_91 : begin
        fsm_output = 8'b01011110;
        state_var_NS = STORE_MAIN_LOOP_C_92;
      end
      STORE_MAIN_LOOP_C_92 : begin
        fsm_output = 8'b01011111;
        state_var_NS = STORE_MAIN_LOOP_C_93;
      end
      STORE_MAIN_LOOP_C_93 : begin
        fsm_output = 8'b01100000;
        state_var_NS = STORE_MAIN_LOOP_C_94;
      end
      STORE_MAIN_LOOP_C_94 : begin
        fsm_output = 8'b01100001;
        state_var_NS = STORE_MAIN_LOOP_C_95;
      end
      STORE_MAIN_LOOP_C_95 : begin
        fsm_output = 8'b01100010;
        state_var_NS = STORE_MAIN_LOOP_C_96;
      end
      STORE_MAIN_LOOP_C_96 : begin
        fsm_output = 8'b01100011;
        state_var_NS = STORE_MAIN_LOOP_C_97;
      end
      STORE_MAIN_LOOP_C_97 : begin
        fsm_output = 8'b01100100;
        state_var_NS = STORE_MAIN_LOOP_C_98;
      end
      STORE_MAIN_LOOP_C_98 : begin
        fsm_output = 8'b01100101;
        state_var_NS = STORE_MAIN_LOOP_C_99;
      end
      STORE_MAIN_LOOP_C_99 : begin
        fsm_output = 8'b01100110;
        state_var_NS = STORE_MAIN_LOOP_C_100;
      end
      STORE_MAIN_LOOP_C_100 : begin
        fsm_output = 8'b01100111;
        state_var_NS = STORE_MAIN_LOOP_C_101;
      end
      STORE_MAIN_LOOP_C_101 : begin
        fsm_output = 8'b01101000;
        state_var_NS = STORE_MAIN_LOOP_C_102;
      end
      STORE_MAIN_LOOP_C_102 : begin
        fsm_output = 8'b01101001;
        state_var_NS = STORE_MAIN_LOOP_C_103;
      end
      STORE_MAIN_LOOP_C_103 : begin
        fsm_output = 8'b01101010;
        state_var_NS = STORE_MAIN_LOOP_C_104;
      end
      STORE_MAIN_LOOP_C_104 : begin
        fsm_output = 8'b01101011;
        state_var_NS = STORE_MAIN_LOOP_C_105;
      end
      STORE_MAIN_LOOP_C_105 : begin
        fsm_output = 8'b01101100;
        state_var_NS = STORE_MAIN_LOOP_C_106;
      end
      STORE_MAIN_LOOP_C_106 : begin
        fsm_output = 8'b01101101;
        state_var_NS = STORE_MAIN_LOOP_C_107;
      end
      STORE_MAIN_LOOP_C_107 : begin
        fsm_output = 8'b01101110;
        state_var_NS = STORE_MAIN_LOOP_C_108;
      end
      STORE_MAIN_LOOP_C_108 : begin
        fsm_output = 8'b01101111;
        state_var_NS = STORE_MAIN_LOOP_C_109;
      end
      STORE_MAIN_LOOP_C_109 : begin
        fsm_output = 8'b01110000;
        state_var_NS = STORE_MAIN_LOOP_C_110;
      end
      STORE_MAIN_LOOP_C_110 : begin
        fsm_output = 8'b01110001;
        state_var_NS = STORE_MAIN_LOOP_C_111;
      end
      STORE_MAIN_LOOP_C_111 : begin
        fsm_output = 8'b01110010;
        state_var_NS = STORE_MAIN_LOOP_C_112;
      end
      STORE_MAIN_LOOP_C_112 : begin
        fsm_output = 8'b01110011;
        state_var_NS = STORE_MAIN_LOOP_C_113;
      end
      STORE_MAIN_LOOP_C_113 : begin
        fsm_output = 8'b01110100;
        state_var_NS = STORE_MAIN_LOOP_C_114;
      end
      STORE_MAIN_LOOP_C_114 : begin
        fsm_output = 8'b01110101;
        state_var_NS = STORE_MAIN_LOOP_C_115;
      end
      STORE_MAIN_LOOP_C_115 : begin
        fsm_output = 8'b01110110;
        state_var_NS = STORE_MAIN_LOOP_C_116;
      end
      STORE_MAIN_LOOP_C_116 : begin
        fsm_output = 8'b01110111;
        state_var_NS = STORE_MAIN_LOOP_C_117;
      end
      STORE_MAIN_LOOP_C_117 : begin
        fsm_output = 8'b01111000;
        state_var_NS = STORE_MAIN_LOOP_C_118;
      end
      STORE_MAIN_LOOP_C_118 : begin
        fsm_output = 8'b01111001;
        state_var_NS = STORE_MAIN_LOOP_C_119;
      end
      STORE_MAIN_LOOP_C_119 : begin
        fsm_output = 8'b01111010;
        state_var_NS = STORE_MAIN_LOOP_C_120;
      end
      STORE_MAIN_LOOP_C_120 : begin
        fsm_output = 8'b01111011;
        state_var_NS = STORE_MAIN_LOOP_C_121;
      end
      STORE_MAIN_LOOP_C_121 : begin
        fsm_output = 8'b01111100;
        state_var_NS = STORE_MAIN_LOOP_C_122;
      end
      STORE_MAIN_LOOP_C_122 : begin
        fsm_output = 8'b01111101;
        state_var_NS = STORE_MAIN_LOOP_C_123;
      end
      STORE_MAIN_LOOP_C_123 : begin
        fsm_output = 8'b01111110;
        state_var_NS = STORE_MAIN_LOOP_C_124;
      end
      STORE_MAIN_LOOP_C_124 : begin
        fsm_output = 8'b01111111;
        state_var_NS = STORE_MAIN_LOOP_C_125;
      end
      STORE_MAIN_LOOP_C_125 : begin
        fsm_output = 8'b10000000;
        state_var_NS = STORE_MAIN_LOOP_C_126;
      end
      STORE_MAIN_LOOP_C_126 : begin
        fsm_output = 8'b10000001;
        state_var_NS = STORE_MAIN_LOOP_C_127;
      end
      STORE_MAIN_LOOP_C_127 : begin
        fsm_output = 8'b10000010;
        state_var_NS = STORE_MAIN_LOOP_C_128;
      end
      STORE_MAIN_LOOP_C_128 : begin
        fsm_output = 8'b10000011;
        state_var_NS = STORE_MAIN_LOOP_C_129;
      end
      STORE_MAIN_LOOP_C_129 : begin
        fsm_output = 8'b10000100;
        state_var_NS = STORE_OUTPUT_INNER_LOOP_C_0;
      end
      STORE_OUTPUT_INNER_LOOP_C_0 : begin
        fsm_output = 8'b10000101;
        if ( STORE_OUTPUT_INNER_LOOP_C_0_tr0 ) begin
          state_var_NS = STORE_MAIN_LOOP_C_130;
        end
        else begin
          state_var_NS = STORE_OUTPUT_INNER_LOOP_C_0;
        end
      end
      STORE_MAIN_LOOP_C_130 : begin
        fsm_output = 8'b10000110;
        if ( STORE_MAIN_LOOP_C_130_tr0 ) begin
          state_var_NS = COMPUTE_BATCH_LOOP_C_1;
        end
        else begin
          state_var_NS = STORE_MAIN_LOOP_C_0;
        end
      end
      COMPUTE_BATCH_LOOP_C_1 : begin
        fsm_output = 8'b10000111;
        if ( COMPUTE_BATCH_LOOP_C_1_tr0 ) begin
          state_var_NS = COMPUTE_BATCH_LOOP_C_0;
        end
        else begin
          state_var_NS = store_output_rlp_C_1;
        end
      end
      store_output_rlp_C_1 : begin
        fsm_output = 8'b10001000;
        state_var_NS = PROCESS_DONE_LOOP_C_0;
      end
      PROCESS_DONE_LOOP_C_0 : begin
        fsm_output = 8'b10001001;
        state_var_NS = PROCESS_DONE_LOOP_C_0;
      end
      // WAIT_FOR_CONFIG_LOOP_C_0
      default : begin
        fsm_output = 8'b00000000;
        if ( WAIT_FOR_CONFIG_LOOP_C_0_tr0 ) begin
          state_var_NS = WAIT_FOR_CONFIG_LOOP_C_0;
        end
        else begin
          state_var_NS = store_output_rlp_C_0;
        end
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= WAIT_FOR_CONFIG_LOOP_C_0;
    end
    else if ( store_output_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_staller
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_staller (
  store_output_wen, output_ready_channel_Push_mioi_wen_comp, dma_write_ctrl_Push_mioi_wen_comp,
      dma_write_chnl_Push_mioi_wen_comp, plm_out_cnsi_wen_comp
);
  output store_output_wen;
  input output_ready_channel_Push_mioi_wen_comp;
  input dma_write_ctrl_Push_mioi_wen_comp;
  input dma_write_chnl_Push_mioi_wen_comp;
  input plm_out_cnsi_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign store_output_wen = output_ready_channel_Push_mioi_wen_comp & dma_write_ctrl_Push_mioi_wen_comp
      & dma_write_chnl_Push_mioi_wen_comp & plm_out_cnsi_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_plm_out_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_plm_out_wait_dp
    (
  clk, rst, plm_out_cnsi_oswt, plm_out_cnsi_wen_comp, plm_out_cnsi_idat_mxwt, plm_out_cnsi_biwt,
      plm_out_cnsi_bdwt, plm_out_cnsi_bcwt, plm_out_cnsi_idat
);
  input clk;
  input rst;
  input plm_out_cnsi_oswt;
  output plm_out_cnsi_wen_comp;
  output [4095:0] plm_out_cnsi_idat_mxwt;
  input plm_out_cnsi_biwt;
  input plm_out_cnsi_bdwt;
  output plm_out_cnsi_bcwt;
  reg plm_out_cnsi_bcwt;
  input [4095:0] plm_out_cnsi_idat;


  // Interconnect Declarations
  reg [4095:0] plm_out_cnsi_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cnsi_wen_comp = (~ plm_out_cnsi_oswt) | plm_out_cnsi_biwt | plm_out_cnsi_bcwt;
  assign plm_out_cnsi_idat_mxwt = MUX_v_4096_2_2(plm_out_cnsi_idat, plm_out_cnsi_idat_bfwt,
      plm_out_cnsi_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cnsi_bcwt <= 1'b0;
    end
    else begin
      plm_out_cnsi_bcwt <= ~((~(plm_out_cnsi_bcwt | plm_out_cnsi_biwt)) | plm_out_cnsi_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( plm_out_cnsi_biwt ) begin
      plm_out_cnsi_idat_bfwt <= plm_out_cnsi_idat;
    end
  end

  function automatic [4095:0] MUX_v_4096_2_2;
    input [4095:0] input_0;
    input [4095:0] input_1;
    input [0:0] sel;
    reg [4095:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4096_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_plm_out_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_plm_out_wait_ctrl
    (
  store_output_wen, plm_out_cnsi_oswt, plm_out_cnsi_biwt, plm_out_cnsi_bdwt, plm_out_cnsi_bcwt,
      plm_out_cnsi_irdy_store_output_sct, plm_out_cnsi_ivld
);
  input store_output_wen;
  input plm_out_cnsi_oswt;
  output plm_out_cnsi_biwt;
  output plm_out_cnsi_bdwt;
  input plm_out_cnsi_bcwt;
  output plm_out_cnsi_irdy_store_output_sct;
  input plm_out_cnsi_ivld;


  // Interconnect Declarations
  wire plm_out_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cnsi_bdwt = plm_out_cnsi_oswt & store_output_wen;
  assign plm_out_cnsi_biwt = plm_out_cnsi_ogwt & plm_out_cnsi_ivld;
  assign plm_out_cnsi_ogwt = plm_out_cnsi_oswt & (~ plm_out_cnsi_bcwt);
  assign plm_out_cnsi_irdy_store_output_sct = plm_out_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp
    (
  clk, rst, dma_write_chnl_Push_mioi_oswt, dma_write_chnl_Push_mioi_wen_comp, dma_write_chnl_Push_mioi_m_rsc_dat_store_output,
      dma_write_chnl_Push_mioi_m_rsc_dat, dma_write_chnl_Push_mioi_biwt, dma_write_chnl_Push_mioi_bdwt,
      dma_write_chnl_Push_mioi_bcwt, dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
);
  input clk;
  input rst;
  input dma_write_chnl_Push_mioi_oswt;
  output dma_write_chnl_Push_mioi_wen_comp;
  input [63:0] dma_write_chnl_Push_mioi_m_rsc_dat_store_output;
  output [63:0] dma_write_chnl_Push_mioi_m_rsc_dat;
  input dma_write_chnl_Push_mioi_biwt;
  input dma_write_chnl_Push_mioi_bdwt;
  output dma_write_chnl_Push_mioi_bcwt;
  reg dma_write_chnl_Push_mioi_bcwt;
  input dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dma_write_chnl_Push_mioi_wen_comp = (~ dma_write_chnl_Push_mioi_oswt) |
      dma_write_chnl_Push_mioi_biwt | dma_write_chnl_Push_mioi_bcwt;
  assign dma_write_chnl_Push_mioi_m_rsc_dat = {dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff)
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff) , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff) , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff) , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff)
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff) , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff) , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , (~ dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff) , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff
      , dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff , (dma_write_chnl_Push_mioi_m_rsc_dat_store_output[31:0])};
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_chnl_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_write_chnl_Push_mioi_bcwt <= ~((~(dma_write_chnl_Push_mioi_bcwt | dma_write_chnl_Push_mioi_biwt))
          | dma_write_chnl_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl
    (
  store_output_wen, dma_write_chnl_Push_mioi_oswt, dma_write_chnl_Push_mioi_biwt,
      dma_write_chnl_Push_mioi_bdwt, dma_write_chnl_Push_mioi_bcwt, dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld,
      dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff, dma_write_chnl_Push_mioi_oswt_pff
);
  input store_output_wen;
  input dma_write_chnl_Push_mioi_oswt;
  output dma_write_chnl_Push_mioi_biwt;
  output dma_write_chnl_Push_mioi_bdwt;
  input dma_write_chnl_Push_mioi_bcwt;
  input dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld;
  output dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff;
  input dma_write_chnl_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dma_write_chnl_Push_mioi_bdwt = dma_write_chnl_Push_mioi_oswt & store_output_wen;
  assign dma_write_chnl_Push_mioi_biwt = dma_write_chnl_Push_mioi_oswt & (~ dma_write_chnl_Push_mioi_bcwt)
      & dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld;
  assign dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff = dma_write_chnl_Push_mioi_oswt_pff
      & store_output_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp
    (
  clk, rst, dma_write_ctrl_Push_mioi_oswt, dma_write_ctrl_Push_mioi_wen_comp, dma_write_ctrl_Push_mioi_biwt,
      dma_write_ctrl_Push_mioi_bdwt, dma_write_ctrl_Push_mioi_bcwt
);
  input clk;
  input rst;
  input dma_write_ctrl_Push_mioi_oswt;
  output dma_write_ctrl_Push_mioi_wen_comp;
  input dma_write_ctrl_Push_mioi_biwt;
  input dma_write_ctrl_Push_mioi_bdwt;
  output dma_write_ctrl_Push_mioi_bcwt;
  reg dma_write_ctrl_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dma_write_ctrl_Push_mioi_wen_comp = (~ dma_write_ctrl_Push_mioi_oswt) |
      dma_write_ctrl_Push_mioi_biwt | dma_write_ctrl_Push_mioi_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_ctrl_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_write_ctrl_Push_mioi_bcwt <= ~((~(dma_write_ctrl_Push_mioi_bcwt | dma_write_ctrl_Push_mioi_biwt))
          | dma_write_ctrl_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl
    (
  store_output_wen, dma_write_ctrl_Push_mioi_oswt, dma_write_ctrl_Push_mioi_biwt,
      dma_write_ctrl_Push_mioi_bdwt, dma_write_ctrl_Push_mioi_bcwt, dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_output_sct,
      dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld, dma_write_ctrl_Push_mioi_oswt_pff
);
  input store_output_wen;
  input dma_write_ctrl_Push_mioi_oswt;
  output dma_write_ctrl_Push_mioi_biwt;
  output dma_write_ctrl_Push_mioi_bdwt;
  input dma_write_ctrl_Push_mioi_bcwt;
  output dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_output_sct;
  input dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  input dma_write_ctrl_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dma_write_ctrl_Push_mioi_bdwt = dma_write_ctrl_Push_mioi_oswt & store_output_wen;
  assign dma_write_ctrl_Push_mioi_biwt = dma_write_ctrl_Push_mioi_oswt & (~ dma_write_ctrl_Push_mioi_bcwt)
      & dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  assign dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_output_sct = dma_write_ctrl_Push_mioi_oswt_pff
      & store_output_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_output_ready_channel_Push_mioi_output_ready_channel_Push_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_output_ready_channel_Push_mioi_output_ready_channel_Push_mio_wait_dp
    (
  clk, rst, output_ready_channel_Push_mioi_oswt, output_ready_channel_Push_mioi_wen_comp,
      output_ready_channel_Push_mioi_biwt, output_ready_channel_Push_mioi_bdwt, output_ready_channel_Push_mioi_bcwt
);
  input clk;
  input rst;
  input output_ready_channel_Push_mioi_oswt;
  output output_ready_channel_Push_mioi_wen_comp;
  input output_ready_channel_Push_mioi_biwt;
  input output_ready_channel_Push_mioi_bdwt;
  output output_ready_channel_Push_mioi_bcwt;
  reg output_ready_channel_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign output_ready_channel_Push_mioi_wen_comp = (~ output_ready_channel_Push_mioi_oswt)
      | output_ready_channel_Push_mioi_biwt | output_ready_channel_Push_mioi_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      output_ready_channel_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      output_ready_channel_Push_mioi_bcwt <= ~((~(output_ready_channel_Push_mioi_bcwt
          | output_ready_channel_Push_mioi_biwt)) | output_ready_channel_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_output_ready_channel_Push_mioi_output_ready_channel_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_output_ready_channel_Push_mioi_output_ready_channel_Push_mio_wait_ctrl
    (
  store_output_wen, output_ready_channel_Push_mioi_oswt, output_ready_channel_Push_mioi_biwt,
      output_ready_channel_Push_mioi_bdwt, output_ready_channel_Push_mioi_bcwt, output_ready_channel_Push_mioi_ccs_ccore_start_rsc_dat_store_output_sct,
      output_ready_channel_Push_mioi_ccs_ccore_done_sync_vld, output_ready_channel_Push_mioi_oswt_pff
);
  input store_output_wen;
  input output_ready_channel_Push_mioi_oswt;
  output output_ready_channel_Push_mioi_biwt;
  output output_ready_channel_Push_mioi_bdwt;
  input output_ready_channel_Push_mioi_bcwt;
  output output_ready_channel_Push_mioi_ccs_ccore_start_rsc_dat_store_output_sct;
  input output_ready_channel_Push_mioi_ccs_ccore_done_sync_vld;
  input output_ready_channel_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign output_ready_channel_Push_mioi_bdwt = output_ready_channel_Push_mioi_oswt
      & store_output_wen;
  assign output_ready_channel_Push_mioi_biwt = output_ready_channel_Push_mioi_oswt
      & (~ output_ready_channel_Push_mioi_bcwt) & output_ready_channel_Push_mioi_ccs_ccore_done_sync_vld;
  assign output_ready_channel_Push_mioi_ccs_ccore_start_rsc_dat_store_output_sct
      = output_ready_channel_Push_mioi_oswt_pff & store_output_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_51_1_1024_2_2_1024_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_51_1_1024_2_2_1024_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [1023:0] qb;
  output web;
  output [1023:0] db;
  output adrb;
  input [1023:0] qa;
  output wea;
  output [1023:0] da;
  output adra;
  input [1:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [2047:0] da_d;
  output [2047:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[2047:1024] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[2047:1024]);
  assign adrb = (adra_d[1]);
  assign qa_d[1023:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[1023:0]);
  assign adra = (adra_d[0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_50_1_1024_2_2_1024_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_50_1_1024_2_2_1024_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [1023:0] qb;
  output web;
  output [1023:0] db;
  output adrb;
  input [1023:0] qa;
  output wea;
  output [1023:0] da;
  output adra;
  input [1:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [2047:0] da_d;
  output [2047:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[2047:1024] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[2047:1024]);
  assign adrb = (adra_d[1]);
  assign qa_d[1023:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[1023:0]);
  assign adra = (adra_d[0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_49_1_1024_2_2_1024_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_49_1_1024_2_2_1024_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [1023:0] qb;
  output web;
  output [1023:0] db;
  output adrb;
  input [1023:0] qa;
  output wea;
  output [1023:0] da;
  output adra;
  input [1:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [2047:0] da_d;
  output [2047:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[2047:1024] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[2047:1024]);
  assign adrb = (adra_d[1]);
  assign qa_d[1023:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[1023:0]);
  assign adra = (adra_d[0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_48_1_1024_2_2_1024_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_48_1_1024_2_2_1024_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [1023:0] qb;
  output web;
  output [1023:0] db;
  output adrb;
  input [1023:0] qa;
  output wea;
  output [1023:0] da;
  output adra;
  input [1:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [2047:0] da_d;
  output [2047:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[2047:1024] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[2047:1024]);
  assign adrb = (adra_d[1]);
  assign qa_d[1023:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[1023:0]);
  assign adra = (adra_d[0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_19_7_67_128_128_67_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_19_7_67_128_128_67_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [66:0] q;
  output [6:0] radr;
  output we;
  output [66:0] d;
  output [6:0] wadr;
  input clken_d;
  input [66:0] d_d;
  output [66:0] q_d;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_compute_kernel_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_compute_kernel_fsm (
  clk, rst, compute_kernel_wen, fsm_output, WAIT_FOR_CONFIG_LOOP_C_0_tr0, compute_kernel_rlp_C_0_tr0,
      COMPUTE_OUTER_LOOP_C_1_tr0, COMPUTE_BATCH_LOOP_C_0_tr0
);
  input clk;
  input rst;
  input compute_kernel_wen;
  output [5:0] fsm_output;
  reg [5:0] fsm_output;
  input WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  input compute_kernel_rlp_C_0_tr0;
  input COMPUTE_OUTER_LOOP_C_1_tr0;
  input COMPUTE_BATCH_LOOP_C_0_tr0;


  // FSM State Type Declaration for esp_acc_softmax_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_1
  parameter
    WAIT_FOR_CONFIG_LOOP_C_0 = 3'd0,
    compute_kernel_rlp_C_0 = 3'd1,
    COMPUTE_OUTER_LOOP_C_0 = 3'd2,
    COMPUTE_OUTER_LOOP_C_1 = 3'd3,
    COMPUTE_BATCH_LOOP_C_0 = 3'd4,
    PROCESS_DONE_LOOP_C_0 = 3'd5;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_softmax_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_1
    case (state_var)
      compute_kernel_rlp_C_0 : begin
        fsm_output = 6'b000010;
        if ( compute_kernel_rlp_C_0_tr0 ) begin
          state_var_NS = COMPUTE_OUTER_LOOP_C_0;
        end
        else begin
          state_var_NS = PROCESS_DONE_LOOP_C_0;
        end
      end
      COMPUTE_OUTER_LOOP_C_0 : begin
        fsm_output = 6'b000100;
        state_var_NS = COMPUTE_OUTER_LOOP_C_1;
      end
      COMPUTE_OUTER_LOOP_C_1 : begin
        fsm_output = 6'b001000;
        if ( COMPUTE_OUTER_LOOP_C_1_tr0 ) begin
          state_var_NS = COMPUTE_OUTER_LOOP_C_0;
        end
        else begin
          state_var_NS = COMPUTE_BATCH_LOOP_C_0;
        end
      end
      COMPUTE_BATCH_LOOP_C_0 : begin
        fsm_output = 6'b010000;
        if ( COMPUTE_BATCH_LOOP_C_0_tr0 ) begin
          state_var_NS = COMPUTE_OUTER_LOOP_C_0;
        end
        else begin
          state_var_NS = PROCESS_DONE_LOOP_C_0;
        end
      end
      PROCESS_DONE_LOOP_C_0 : begin
        fsm_output = 6'b100000;
        state_var_NS = PROCESS_DONE_LOOP_C_0;
      end
      // WAIT_FOR_CONFIG_LOOP_C_0
      default : begin
        fsm_output = 6'b000001;
        if ( WAIT_FOR_CONFIG_LOOP_C_0_tr0 ) begin
          state_var_NS = WAIT_FOR_CONFIG_LOOP_C_0;
        end
        else begin
          state_var_NS = compute_kernel_rlp_C_0;
        end
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= WAIT_FOR_CONFIG_LOOP_C_0;
    end
    else if ( compute_kernel_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_staller
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_staller (
  compute_kernel_wen, input_ready_channel_Push_mioi_wen_comp, output_ready_channel_Pop_mioi_wen_comp,
      plm_in_cnsi_wen_comp, plm_out_cnsi_wen_comp
);
  output compute_kernel_wen;
  input input_ready_channel_Push_mioi_wen_comp;
  input output_ready_channel_Pop_mioi_wen_comp;
  input plm_in_cnsi_wen_comp;
  input plm_out_cnsi_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign compute_kernel_wen = input_ready_channel_Push_mioi_wen_comp & output_ready_channel_Pop_mioi_wen_comp
      & plm_in_cnsi_wen_comp & plm_out_cnsi_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi_plm_out_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi_plm_out_wait_dp
    (
  clk, rst, plm_out_cnsi_oswt, plm_out_cnsi_wen_comp, plm_out_cnsi_biwt, plm_out_cnsi_bdwt,
      plm_out_cnsi_bcwt
);
  input clk;
  input rst;
  input plm_out_cnsi_oswt;
  output plm_out_cnsi_wen_comp;
  input plm_out_cnsi_biwt;
  input plm_out_cnsi_bdwt;
  output plm_out_cnsi_bcwt;
  reg plm_out_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cnsi_wen_comp = (~ plm_out_cnsi_oswt) | plm_out_cnsi_biwt | plm_out_cnsi_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_out_cnsi_bcwt <= 1'b0;
    end
    else begin
      plm_out_cnsi_bcwt <= ~((~(plm_out_cnsi_bcwt | plm_out_cnsi_biwt)) | plm_out_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi_plm_out_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi_plm_out_wait_ctrl
    (
  compute_kernel_wen, plm_out_cnsi_oswt, plm_out_cnsi_irdy, plm_out_cnsi_biwt, plm_out_cnsi_bdwt,
      plm_out_cnsi_bcwt, plm_out_cnsi_ivld_compute_kernel_sct
);
  input compute_kernel_wen;
  input plm_out_cnsi_oswt;
  input plm_out_cnsi_irdy;
  output plm_out_cnsi_biwt;
  output plm_out_cnsi_bdwt;
  input plm_out_cnsi_bcwt;
  output plm_out_cnsi_ivld_compute_kernel_sct;


  // Interconnect Declarations
  wire plm_out_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_out_cnsi_bdwt = plm_out_cnsi_oswt & compute_kernel_wen;
  assign plm_out_cnsi_biwt = plm_out_cnsi_ogwt & plm_out_cnsi_irdy;
  assign plm_out_cnsi_ogwt = plm_out_cnsi_oswt & (~ plm_out_cnsi_bcwt);
  assign plm_out_cnsi_ivld_compute_kernel_sct = plm_out_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_plm_in_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_plm_in_wait_dp
    (
  clk, rst, plm_in_cnsi_oswt, plm_in_cnsi_wen_comp, plm_in_cnsi_idat_mxwt, plm_in_cnsi_biwt,
      plm_in_cnsi_bdwt, plm_in_cnsi_bcwt, plm_in_cnsi_idat
);
  input clk;
  input rst;
  input plm_in_cnsi_oswt;
  output plm_in_cnsi_wen_comp;
  output [4095:0] plm_in_cnsi_idat_mxwt;
  input plm_in_cnsi_biwt;
  input plm_in_cnsi_bdwt;
  output plm_in_cnsi_bcwt;
  reg plm_in_cnsi_bcwt;
  input [4095:0] plm_in_cnsi_idat;


  // Interconnect Declarations
  reg [4095:0] plm_in_cnsi_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cnsi_wen_comp = (~ plm_in_cnsi_oswt) | plm_in_cnsi_biwt | plm_in_cnsi_bcwt;
  assign plm_in_cnsi_idat_mxwt = MUX_v_4096_2_2(plm_in_cnsi_idat, plm_in_cnsi_idat_bfwt,
      plm_in_cnsi_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cnsi_bcwt <= 1'b0;
    end
    else begin
      plm_in_cnsi_bcwt <= ~((~(plm_in_cnsi_bcwt | plm_in_cnsi_biwt)) | plm_in_cnsi_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( plm_in_cnsi_biwt ) begin
      plm_in_cnsi_idat_bfwt <= plm_in_cnsi_idat;
    end
  end

  function automatic [4095:0] MUX_v_4096_2_2;
    input [4095:0] input_0;
    input [4095:0] input_1;
    input [0:0] sel;
    reg [4095:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4096_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_plm_in_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_plm_in_wait_ctrl
    (
  compute_kernel_wen, plm_in_cnsi_oswt, plm_in_cnsi_biwt, plm_in_cnsi_bdwt, plm_in_cnsi_bcwt,
      plm_in_cnsi_irdy_compute_kernel_sct, plm_in_cnsi_ivld
);
  input compute_kernel_wen;
  input plm_in_cnsi_oswt;
  output plm_in_cnsi_biwt;
  output plm_in_cnsi_bdwt;
  input plm_in_cnsi_bcwt;
  output plm_in_cnsi_irdy_compute_kernel_sct;
  input plm_in_cnsi_ivld;


  // Interconnect Declarations
  wire plm_in_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cnsi_bdwt = plm_in_cnsi_oswt & compute_kernel_wen;
  assign plm_in_cnsi_biwt = plm_in_cnsi_ogwt & plm_in_cnsi_ivld;
  assign plm_in_cnsi_ogwt = plm_in_cnsi_oswt & (~ plm_in_cnsi_bcwt);
  assign plm_in_cnsi_irdy_compute_kernel_sct = plm_in_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_channel_Pop_mioi_output_ready_channel_Pop_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_channel_Pop_mioi_output_ready_channel_Pop_mio_wait_dp
    (
  clk, rst, output_ready_channel_Pop_mioi_oswt, output_ready_channel_Pop_mioi_wen_comp,
      output_ready_channel_Pop_mioi_biwt, output_ready_channel_Pop_mioi_bdwt, output_ready_channel_Pop_mioi_bcwt
);
  input clk;
  input rst;
  input output_ready_channel_Pop_mioi_oswt;
  output output_ready_channel_Pop_mioi_wen_comp;
  input output_ready_channel_Pop_mioi_biwt;
  input output_ready_channel_Pop_mioi_bdwt;
  output output_ready_channel_Pop_mioi_bcwt;
  reg output_ready_channel_Pop_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign output_ready_channel_Pop_mioi_wen_comp = (~ output_ready_channel_Pop_mioi_oswt)
      | output_ready_channel_Pop_mioi_biwt | output_ready_channel_Pop_mioi_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      output_ready_channel_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      output_ready_channel_Pop_mioi_bcwt <= ~((~(output_ready_channel_Pop_mioi_bcwt
          | output_ready_channel_Pop_mioi_biwt)) | output_ready_channel_Pop_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_channel_Pop_mioi_output_ready_channel_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_channel_Pop_mioi_output_ready_channel_Pop_mio_wait_ctrl
    (
  compute_kernel_wen, output_ready_channel_Pop_mioi_oswt, output_ready_channel_Pop_mioi_biwt,
      output_ready_channel_Pop_mioi_bdwt, output_ready_channel_Pop_mioi_bcwt, output_ready_channel_Pop_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct,
      output_ready_channel_Pop_mioi_ccs_ccore_done_sync_vld, output_ready_channel_Pop_mioi_oswt_pff
);
  input compute_kernel_wen;
  input output_ready_channel_Pop_mioi_oswt;
  output output_ready_channel_Pop_mioi_biwt;
  output output_ready_channel_Pop_mioi_bdwt;
  input output_ready_channel_Pop_mioi_bcwt;
  output output_ready_channel_Pop_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct;
  input output_ready_channel_Pop_mioi_ccs_ccore_done_sync_vld;
  input output_ready_channel_Pop_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign output_ready_channel_Pop_mioi_bdwt = output_ready_channel_Pop_mioi_oswt
      & compute_kernel_wen;
  assign output_ready_channel_Pop_mioi_biwt = output_ready_channel_Pop_mioi_oswt
      & (~ output_ready_channel_Pop_mioi_bcwt) & output_ready_channel_Pop_mioi_ccs_ccore_done_sync_vld;
  assign output_ready_channel_Pop_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct
      = output_ready_channel_Pop_mioi_oswt_pff & compute_kernel_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_channel_Push_mioi_input_ready_channel_Push_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_channel_Push_mioi_input_ready_channel_Push_mio_wait_dp
    (
  clk, rst, input_ready_channel_Push_mioi_oswt, input_ready_channel_Push_mioi_wen_comp,
      input_ready_channel_Push_mioi_biwt, input_ready_channel_Push_mioi_bdwt, input_ready_channel_Push_mioi_bcwt
);
  input clk;
  input rst;
  input input_ready_channel_Push_mioi_oswt;
  output input_ready_channel_Push_mioi_wen_comp;
  input input_ready_channel_Push_mioi_biwt;
  input input_ready_channel_Push_mioi_bdwt;
  output input_ready_channel_Push_mioi_bcwt;
  reg input_ready_channel_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign input_ready_channel_Push_mioi_wen_comp = (~ input_ready_channel_Push_mioi_oswt)
      | input_ready_channel_Push_mioi_biwt | input_ready_channel_Push_mioi_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      input_ready_channel_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      input_ready_channel_Push_mioi_bcwt <= ~((~(input_ready_channel_Push_mioi_bcwt
          | input_ready_channel_Push_mioi_biwt)) | input_ready_channel_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_channel_Push_mioi_input_ready_channel_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_channel_Push_mioi_input_ready_channel_Push_mio_wait_ctrl
    (
  compute_kernel_wen, input_ready_channel_Push_mioi_oswt, input_ready_channel_Push_mioi_biwt,
      input_ready_channel_Push_mioi_bdwt, input_ready_channel_Push_mioi_bcwt, input_ready_channel_Push_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct,
      input_ready_channel_Push_mioi_ccs_ccore_done_sync_vld, input_ready_channel_Push_mioi_oswt_pff
);
  input compute_kernel_wen;
  input input_ready_channel_Push_mioi_oswt;
  output input_ready_channel_Push_mioi_biwt;
  output input_ready_channel_Push_mioi_bdwt;
  input input_ready_channel_Push_mioi_bcwt;
  output input_ready_channel_Push_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct;
  input input_ready_channel_Push_mioi_ccs_ccore_done_sync_vld;
  input input_ready_channel_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign input_ready_channel_Push_mioi_bdwt = input_ready_channel_Push_mioi_oswt
      & compute_kernel_wen;
  assign input_ready_channel_Push_mioi_biwt = input_ready_channel_Push_mioi_oswt
      & (~ input_ready_channel_Push_mioi_bcwt) & input_ready_channel_Push_mioi_ccs_ccore_done_sync_vld;
  assign input_ready_channel_Push_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct
      = input_ready_channel_Push_mioi_oswt_pff & compute_kernel_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_16_7_32_128_128_32_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_16_7_32_128_128_32_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [31:0] q;
  output [6:0] radr;
  output we;
  output [31:0] d;
  output [6:0] wadr;
  input clken_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_load_input_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_load_input_fsm (
  clk, rst, load_input_wen, fsm_output, WAIT_FOR_CONFIG_LOOP_C_0_tr0, load_input_rlp_C_0_tr0,
      LOAD_BATCH_LOOP_C_0_tr0, LOAD_DATA_INNER_LOOP_C_0_tr0, LOAD_DATA_OUTER_LOOP_C_131_tr0,
      LOAD_BATCH_LOOP_C_1_tr0
);
  input clk;
  input rst;
  input load_input_wen;
  output [7:0] fsm_output;
  reg [7:0] fsm_output;
  input WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  input load_input_rlp_C_0_tr0;
  input LOAD_BATCH_LOOP_C_0_tr0;
  input LOAD_DATA_INNER_LOOP_C_0_tr0;
  input LOAD_DATA_OUTER_LOOP_C_131_tr0;
  input LOAD_BATCH_LOOP_C_1_tr0;


  // FSM State Type Declaration for esp_acc_softmax_softmax_load_input_load_input_load_input_fsm_1
  parameter
    WAIT_FOR_CONFIG_LOOP_C_0 = 8'd0,
    load_input_rlp_C_0 = 8'd1,
    LOAD_BATCH_LOOP_C_0 = 8'd2,
    LOAD_DATA_OUTER_LOOP_C_0 = 8'd3,
    LOAD_DATA_OUTER_LOOP_C_1 = 8'd4,
    LOAD_DATA_INNER_LOOP_C_0 = 8'd5,
    LOAD_DATA_OUTER_LOOP_C_2 = 8'd6,
    LOAD_DATA_OUTER_LOOP_C_3 = 8'd7,
    LOAD_DATA_OUTER_LOOP_C_4 = 8'd8,
    LOAD_DATA_OUTER_LOOP_C_5 = 8'd9,
    LOAD_DATA_OUTER_LOOP_C_6 = 8'd10,
    LOAD_DATA_OUTER_LOOP_C_7 = 8'd11,
    LOAD_DATA_OUTER_LOOP_C_8 = 8'd12,
    LOAD_DATA_OUTER_LOOP_C_9 = 8'd13,
    LOAD_DATA_OUTER_LOOP_C_10 = 8'd14,
    LOAD_DATA_OUTER_LOOP_C_11 = 8'd15,
    LOAD_DATA_OUTER_LOOP_C_12 = 8'd16,
    LOAD_DATA_OUTER_LOOP_C_13 = 8'd17,
    LOAD_DATA_OUTER_LOOP_C_14 = 8'd18,
    LOAD_DATA_OUTER_LOOP_C_15 = 8'd19,
    LOAD_DATA_OUTER_LOOP_C_16 = 8'd20,
    LOAD_DATA_OUTER_LOOP_C_17 = 8'd21,
    LOAD_DATA_OUTER_LOOP_C_18 = 8'd22,
    LOAD_DATA_OUTER_LOOP_C_19 = 8'd23,
    LOAD_DATA_OUTER_LOOP_C_20 = 8'd24,
    LOAD_DATA_OUTER_LOOP_C_21 = 8'd25,
    LOAD_DATA_OUTER_LOOP_C_22 = 8'd26,
    LOAD_DATA_OUTER_LOOP_C_23 = 8'd27,
    LOAD_DATA_OUTER_LOOP_C_24 = 8'd28,
    LOAD_DATA_OUTER_LOOP_C_25 = 8'd29,
    LOAD_DATA_OUTER_LOOP_C_26 = 8'd30,
    LOAD_DATA_OUTER_LOOP_C_27 = 8'd31,
    LOAD_DATA_OUTER_LOOP_C_28 = 8'd32,
    LOAD_DATA_OUTER_LOOP_C_29 = 8'd33,
    LOAD_DATA_OUTER_LOOP_C_30 = 8'd34,
    LOAD_DATA_OUTER_LOOP_C_31 = 8'd35,
    LOAD_DATA_OUTER_LOOP_C_32 = 8'd36,
    LOAD_DATA_OUTER_LOOP_C_33 = 8'd37,
    LOAD_DATA_OUTER_LOOP_C_34 = 8'd38,
    LOAD_DATA_OUTER_LOOP_C_35 = 8'd39,
    LOAD_DATA_OUTER_LOOP_C_36 = 8'd40,
    LOAD_DATA_OUTER_LOOP_C_37 = 8'd41,
    LOAD_DATA_OUTER_LOOP_C_38 = 8'd42,
    LOAD_DATA_OUTER_LOOP_C_39 = 8'd43,
    LOAD_DATA_OUTER_LOOP_C_40 = 8'd44,
    LOAD_DATA_OUTER_LOOP_C_41 = 8'd45,
    LOAD_DATA_OUTER_LOOP_C_42 = 8'd46,
    LOAD_DATA_OUTER_LOOP_C_43 = 8'd47,
    LOAD_DATA_OUTER_LOOP_C_44 = 8'd48,
    LOAD_DATA_OUTER_LOOP_C_45 = 8'd49,
    LOAD_DATA_OUTER_LOOP_C_46 = 8'd50,
    LOAD_DATA_OUTER_LOOP_C_47 = 8'd51,
    LOAD_DATA_OUTER_LOOP_C_48 = 8'd52,
    LOAD_DATA_OUTER_LOOP_C_49 = 8'd53,
    LOAD_DATA_OUTER_LOOP_C_50 = 8'd54,
    LOAD_DATA_OUTER_LOOP_C_51 = 8'd55,
    LOAD_DATA_OUTER_LOOP_C_52 = 8'd56,
    LOAD_DATA_OUTER_LOOP_C_53 = 8'd57,
    LOAD_DATA_OUTER_LOOP_C_54 = 8'd58,
    LOAD_DATA_OUTER_LOOP_C_55 = 8'd59,
    LOAD_DATA_OUTER_LOOP_C_56 = 8'd60,
    LOAD_DATA_OUTER_LOOP_C_57 = 8'd61,
    LOAD_DATA_OUTER_LOOP_C_58 = 8'd62,
    LOAD_DATA_OUTER_LOOP_C_59 = 8'd63,
    LOAD_DATA_OUTER_LOOP_C_60 = 8'd64,
    LOAD_DATA_OUTER_LOOP_C_61 = 8'd65,
    LOAD_DATA_OUTER_LOOP_C_62 = 8'd66,
    LOAD_DATA_OUTER_LOOP_C_63 = 8'd67,
    LOAD_DATA_OUTER_LOOP_C_64 = 8'd68,
    LOAD_DATA_OUTER_LOOP_C_65 = 8'd69,
    LOAD_DATA_OUTER_LOOP_C_66 = 8'd70,
    LOAD_DATA_OUTER_LOOP_C_67 = 8'd71,
    LOAD_DATA_OUTER_LOOP_C_68 = 8'd72,
    LOAD_DATA_OUTER_LOOP_C_69 = 8'd73,
    LOAD_DATA_OUTER_LOOP_C_70 = 8'd74,
    LOAD_DATA_OUTER_LOOP_C_71 = 8'd75,
    LOAD_DATA_OUTER_LOOP_C_72 = 8'd76,
    LOAD_DATA_OUTER_LOOP_C_73 = 8'd77,
    LOAD_DATA_OUTER_LOOP_C_74 = 8'd78,
    LOAD_DATA_OUTER_LOOP_C_75 = 8'd79,
    LOAD_DATA_OUTER_LOOP_C_76 = 8'd80,
    LOAD_DATA_OUTER_LOOP_C_77 = 8'd81,
    LOAD_DATA_OUTER_LOOP_C_78 = 8'd82,
    LOAD_DATA_OUTER_LOOP_C_79 = 8'd83,
    LOAD_DATA_OUTER_LOOP_C_80 = 8'd84,
    LOAD_DATA_OUTER_LOOP_C_81 = 8'd85,
    LOAD_DATA_OUTER_LOOP_C_82 = 8'd86,
    LOAD_DATA_OUTER_LOOP_C_83 = 8'd87,
    LOAD_DATA_OUTER_LOOP_C_84 = 8'd88,
    LOAD_DATA_OUTER_LOOP_C_85 = 8'd89,
    LOAD_DATA_OUTER_LOOP_C_86 = 8'd90,
    LOAD_DATA_OUTER_LOOP_C_87 = 8'd91,
    LOAD_DATA_OUTER_LOOP_C_88 = 8'd92,
    LOAD_DATA_OUTER_LOOP_C_89 = 8'd93,
    LOAD_DATA_OUTER_LOOP_C_90 = 8'd94,
    LOAD_DATA_OUTER_LOOP_C_91 = 8'd95,
    LOAD_DATA_OUTER_LOOP_C_92 = 8'd96,
    LOAD_DATA_OUTER_LOOP_C_93 = 8'd97,
    LOAD_DATA_OUTER_LOOP_C_94 = 8'd98,
    LOAD_DATA_OUTER_LOOP_C_95 = 8'd99,
    LOAD_DATA_OUTER_LOOP_C_96 = 8'd100,
    LOAD_DATA_OUTER_LOOP_C_97 = 8'd101,
    LOAD_DATA_OUTER_LOOP_C_98 = 8'd102,
    LOAD_DATA_OUTER_LOOP_C_99 = 8'd103,
    LOAD_DATA_OUTER_LOOP_C_100 = 8'd104,
    LOAD_DATA_OUTER_LOOP_C_101 = 8'd105,
    LOAD_DATA_OUTER_LOOP_C_102 = 8'd106,
    LOAD_DATA_OUTER_LOOP_C_103 = 8'd107,
    LOAD_DATA_OUTER_LOOP_C_104 = 8'd108,
    LOAD_DATA_OUTER_LOOP_C_105 = 8'd109,
    LOAD_DATA_OUTER_LOOP_C_106 = 8'd110,
    LOAD_DATA_OUTER_LOOP_C_107 = 8'd111,
    LOAD_DATA_OUTER_LOOP_C_108 = 8'd112,
    LOAD_DATA_OUTER_LOOP_C_109 = 8'd113,
    LOAD_DATA_OUTER_LOOP_C_110 = 8'd114,
    LOAD_DATA_OUTER_LOOP_C_111 = 8'd115,
    LOAD_DATA_OUTER_LOOP_C_112 = 8'd116,
    LOAD_DATA_OUTER_LOOP_C_113 = 8'd117,
    LOAD_DATA_OUTER_LOOP_C_114 = 8'd118,
    LOAD_DATA_OUTER_LOOP_C_115 = 8'd119,
    LOAD_DATA_OUTER_LOOP_C_116 = 8'd120,
    LOAD_DATA_OUTER_LOOP_C_117 = 8'd121,
    LOAD_DATA_OUTER_LOOP_C_118 = 8'd122,
    LOAD_DATA_OUTER_LOOP_C_119 = 8'd123,
    LOAD_DATA_OUTER_LOOP_C_120 = 8'd124,
    LOAD_DATA_OUTER_LOOP_C_121 = 8'd125,
    LOAD_DATA_OUTER_LOOP_C_122 = 8'd126,
    LOAD_DATA_OUTER_LOOP_C_123 = 8'd127,
    LOAD_DATA_OUTER_LOOP_C_124 = 8'd128,
    LOAD_DATA_OUTER_LOOP_C_125 = 8'd129,
    LOAD_DATA_OUTER_LOOP_C_126 = 8'd130,
    LOAD_DATA_OUTER_LOOP_C_127 = 8'd131,
    LOAD_DATA_OUTER_LOOP_C_128 = 8'd132,
    LOAD_DATA_OUTER_LOOP_C_129 = 8'd133,
    LOAD_DATA_OUTER_LOOP_C_130 = 8'd134,
    LOAD_DATA_OUTER_LOOP_C_131 = 8'd135,
    LOAD_BATCH_LOOP_C_1 = 8'd136,
    PROCESS_DONE_LOOP_C_0 = 8'd137;

  reg [7:0] state_var;
  reg [7:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_softmax_softmax_load_input_load_input_load_input_fsm_1
    case (state_var)
      load_input_rlp_C_0 : begin
        fsm_output = 8'b00000001;
        if ( load_input_rlp_C_0_tr0 ) begin
          state_var_NS = LOAD_BATCH_LOOP_C_0;
        end
        else begin
          state_var_NS = PROCESS_DONE_LOOP_C_0;
        end
      end
      LOAD_BATCH_LOOP_C_0 : begin
        fsm_output = 8'b00000010;
        if ( LOAD_BATCH_LOOP_C_0_tr0 ) begin
          state_var_NS = LOAD_BATCH_LOOP_C_1;
        end
        else begin
          state_var_NS = LOAD_DATA_OUTER_LOOP_C_0;
        end
      end
      LOAD_DATA_OUTER_LOOP_C_0 : begin
        fsm_output = 8'b00000011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_1;
      end
      LOAD_DATA_OUTER_LOOP_C_1 : begin
        fsm_output = 8'b00000100;
        state_var_NS = LOAD_DATA_INNER_LOOP_C_0;
      end
      LOAD_DATA_INNER_LOOP_C_0 : begin
        fsm_output = 8'b00000101;
        if ( LOAD_DATA_INNER_LOOP_C_0_tr0 ) begin
          state_var_NS = LOAD_DATA_OUTER_LOOP_C_2;
        end
        else begin
          state_var_NS = LOAD_DATA_INNER_LOOP_C_0;
        end
      end
      LOAD_DATA_OUTER_LOOP_C_2 : begin
        fsm_output = 8'b00000110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_3;
      end
      LOAD_DATA_OUTER_LOOP_C_3 : begin
        fsm_output = 8'b00000111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_4;
      end
      LOAD_DATA_OUTER_LOOP_C_4 : begin
        fsm_output = 8'b00001000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_5;
      end
      LOAD_DATA_OUTER_LOOP_C_5 : begin
        fsm_output = 8'b00001001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_6;
      end
      LOAD_DATA_OUTER_LOOP_C_6 : begin
        fsm_output = 8'b00001010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_7;
      end
      LOAD_DATA_OUTER_LOOP_C_7 : begin
        fsm_output = 8'b00001011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_8;
      end
      LOAD_DATA_OUTER_LOOP_C_8 : begin
        fsm_output = 8'b00001100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_9;
      end
      LOAD_DATA_OUTER_LOOP_C_9 : begin
        fsm_output = 8'b00001101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_10;
      end
      LOAD_DATA_OUTER_LOOP_C_10 : begin
        fsm_output = 8'b00001110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_11;
      end
      LOAD_DATA_OUTER_LOOP_C_11 : begin
        fsm_output = 8'b00001111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_12;
      end
      LOAD_DATA_OUTER_LOOP_C_12 : begin
        fsm_output = 8'b00010000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_13;
      end
      LOAD_DATA_OUTER_LOOP_C_13 : begin
        fsm_output = 8'b00010001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_14;
      end
      LOAD_DATA_OUTER_LOOP_C_14 : begin
        fsm_output = 8'b00010010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_15;
      end
      LOAD_DATA_OUTER_LOOP_C_15 : begin
        fsm_output = 8'b00010011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_16;
      end
      LOAD_DATA_OUTER_LOOP_C_16 : begin
        fsm_output = 8'b00010100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_17;
      end
      LOAD_DATA_OUTER_LOOP_C_17 : begin
        fsm_output = 8'b00010101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_18;
      end
      LOAD_DATA_OUTER_LOOP_C_18 : begin
        fsm_output = 8'b00010110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_19;
      end
      LOAD_DATA_OUTER_LOOP_C_19 : begin
        fsm_output = 8'b00010111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_20;
      end
      LOAD_DATA_OUTER_LOOP_C_20 : begin
        fsm_output = 8'b00011000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_21;
      end
      LOAD_DATA_OUTER_LOOP_C_21 : begin
        fsm_output = 8'b00011001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_22;
      end
      LOAD_DATA_OUTER_LOOP_C_22 : begin
        fsm_output = 8'b00011010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_23;
      end
      LOAD_DATA_OUTER_LOOP_C_23 : begin
        fsm_output = 8'b00011011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_24;
      end
      LOAD_DATA_OUTER_LOOP_C_24 : begin
        fsm_output = 8'b00011100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_25;
      end
      LOAD_DATA_OUTER_LOOP_C_25 : begin
        fsm_output = 8'b00011101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_26;
      end
      LOAD_DATA_OUTER_LOOP_C_26 : begin
        fsm_output = 8'b00011110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_27;
      end
      LOAD_DATA_OUTER_LOOP_C_27 : begin
        fsm_output = 8'b00011111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_28;
      end
      LOAD_DATA_OUTER_LOOP_C_28 : begin
        fsm_output = 8'b00100000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_29;
      end
      LOAD_DATA_OUTER_LOOP_C_29 : begin
        fsm_output = 8'b00100001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_30;
      end
      LOAD_DATA_OUTER_LOOP_C_30 : begin
        fsm_output = 8'b00100010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_31;
      end
      LOAD_DATA_OUTER_LOOP_C_31 : begin
        fsm_output = 8'b00100011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_32;
      end
      LOAD_DATA_OUTER_LOOP_C_32 : begin
        fsm_output = 8'b00100100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_33;
      end
      LOAD_DATA_OUTER_LOOP_C_33 : begin
        fsm_output = 8'b00100101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_34;
      end
      LOAD_DATA_OUTER_LOOP_C_34 : begin
        fsm_output = 8'b00100110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_35;
      end
      LOAD_DATA_OUTER_LOOP_C_35 : begin
        fsm_output = 8'b00100111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_36;
      end
      LOAD_DATA_OUTER_LOOP_C_36 : begin
        fsm_output = 8'b00101000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_37;
      end
      LOAD_DATA_OUTER_LOOP_C_37 : begin
        fsm_output = 8'b00101001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_38;
      end
      LOAD_DATA_OUTER_LOOP_C_38 : begin
        fsm_output = 8'b00101010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_39;
      end
      LOAD_DATA_OUTER_LOOP_C_39 : begin
        fsm_output = 8'b00101011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_40;
      end
      LOAD_DATA_OUTER_LOOP_C_40 : begin
        fsm_output = 8'b00101100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_41;
      end
      LOAD_DATA_OUTER_LOOP_C_41 : begin
        fsm_output = 8'b00101101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_42;
      end
      LOAD_DATA_OUTER_LOOP_C_42 : begin
        fsm_output = 8'b00101110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_43;
      end
      LOAD_DATA_OUTER_LOOP_C_43 : begin
        fsm_output = 8'b00101111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_44;
      end
      LOAD_DATA_OUTER_LOOP_C_44 : begin
        fsm_output = 8'b00110000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_45;
      end
      LOAD_DATA_OUTER_LOOP_C_45 : begin
        fsm_output = 8'b00110001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_46;
      end
      LOAD_DATA_OUTER_LOOP_C_46 : begin
        fsm_output = 8'b00110010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_47;
      end
      LOAD_DATA_OUTER_LOOP_C_47 : begin
        fsm_output = 8'b00110011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_48;
      end
      LOAD_DATA_OUTER_LOOP_C_48 : begin
        fsm_output = 8'b00110100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_49;
      end
      LOAD_DATA_OUTER_LOOP_C_49 : begin
        fsm_output = 8'b00110101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_50;
      end
      LOAD_DATA_OUTER_LOOP_C_50 : begin
        fsm_output = 8'b00110110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_51;
      end
      LOAD_DATA_OUTER_LOOP_C_51 : begin
        fsm_output = 8'b00110111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_52;
      end
      LOAD_DATA_OUTER_LOOP_C_52 : begin
        fsm_output = 8'b00111000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_53;
      end
      LOAD_DATA_OUTER_LOOP_C_53 : begin
        fsm_output = 8'b00111001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_54;
      end
      LOAD_DATA_OUTER_LOOP_C_54 : begin
        fsm_output = 8'b00111010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_55;
      end
      LOAD_DATA_OUTER_LOOP_C_55 : begin
        fsm_output = 8'b00111011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_56;
      end
      LOAD_DATA_OUTER_LOOP_C_56 : begin
        fsm_output = 8'b00111100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_57;
      end
      LOAD_DATA_OUTER_LOOP_C_57 : begin
        fsm_output = 8'b00111101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_58;
      end
      LOAD_DATA_OUTER_LOOP_C_58 : begin
        fsm_output = 8'b00111110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_59;
      end
      LOAD_DATA_OUTER_LOOP_C_59 : begin
        fsm_output = 8'b00111111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_60;
      end
      LOAD_DATA_OUTER_LOOP_C_60 : begin
        fsm_output = 8'b01000000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_61;
      end
      LOAD_DATA_OUTER_LOOP_C_61 : begin
        fsm_output = 8'b01000001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_62;
      end
      LOAD_DATA_OUTER_LOOP_C_62 : begin
        fsm_output = 8'b01000010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_63;
      end
      LOAD_DATA_OUTER_LOOP_C_63 : begin
        fsm_output = 8'b01000011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_64;
      end
      LOAD_DATA_OUTER_LOOP_C_64 : begin
        fsm_output = 8'b01000100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_65;
      end
      LOAD_DATA_OUTER_LOOP_C_65 : begin
        fsm_output = 8'b01000101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_66;
      end
      LOAD_DATA_OUTER_LOOP_C_66 : begin
        fsm_output = 8'b01000110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_67;
      end
      LOAD_DATA_OUTER_LOOP_C_67 : begin
        fsm_output = 8'b01000111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_68;
      end
      LOAD_DATA_OUTER_LOOP_C_68 : begin
        fsm_output = 8'b01001000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_69;
      end
      LOAD_DATA_OUTER_LOOP_C_69 : begin
        fsm_output = 8'b01001001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_70;
      end
      LOAD_DATA_OUTER_LOOP_C_70 : begin
        fsm_output = 8'b01001010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_71;
      end
      LOAD_DATA_OUTER_LOOP_C_71 : begin
        fsm_output = 8'b01001011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_72;
      end
      LOAD_DATA_OUTER_LOOP_C_72 : begin
        fsm_output = 8'b01001100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_73;
      end
      LOAD_DATA_OUTER_LOOP_C_73 : begin
        fsm_output = 8'b01001101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_74;
      end
      LOAD_DATA_OUTER_LOOP_C_74 : begin
        fsm_output = 8'b01001110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_75;
      end
      LOAD_DATA_OUTER_LOOP_C_75 : begin
        fsm_output = 8'b01001111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_76;
      end
      LOAD_DATA_OUTER_LOOP_C_76 : begin
        fsm_output = 8'b01010000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_77;
      end
      LOAD_DATA_OUTER_LOOP_C_77 : begin
        fsm_output = 8'b01010001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_78;
      end
      LOAD_DATA_OUTER_LOOP_C_78 : begin
        fsm_output = 8'b01010010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_79;
      end
      LOAD_DATA_OUTER_LOOP_C_79 : begin
        fsm_output = 8'b01010011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_80;
      end
      LOAD_DATA_OUTER_LOOP_C_80 : begin
        fsm_output = 8'b01010100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_81;
      end
      LOAD_DATA_OUTER_LOOP_C_81 : begin
        fsm_output = 8'b01010101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_82;
      end
      LOAD_DATA_OUTER_LOOP_C_82 : begin
        fsm_output = 8'b01010110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_83;
      end
      LOAD_DATA_OUTER_LOOP_C_83 : begin
        fsm_output = 8'b01010111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_84;
      end
      LOAD_DATA_OUTER_LOOP_C_84 : begin
        fsm_output = 8'b01011000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_85;
      end
      LOAD_DATA_OUTER_LOOP_C_85 : begin
        fsm_output = 8'b01011001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_86;
      end
      LOAD_DATA_OUTER_LOOP_C_86 : begin
        fsm_output = 8'b01011010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_87;
      end
      LOAD_DATA_OUTER_LOOP_C_87 : begin
        fsm_output = 8'b01011011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_88;
      end
      LOAD_DATA_OUTER_LOOP_C_88 : begin
        fsm_output = 8'b01011100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_89;
      end
      LOAD_DATA_OUTER_LOOP_C_89 : begin
        fsm_output = 8'b01011101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_90;
      end
      LOAD_DATA_OUTER_LOOP_C_90 : begin
        fsm_output = 8'b01011110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_91;
      end
      LOAD_DATA_OUTER_LOOP_C_91 : begin
        fsm_output = 8'b01011111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_92;
      end
      LOAD_DATA_OUTER_LOOP_C_92 : begin
        fsm_output = 8'b01100000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_93;
      end
      LOAD_DATA_OUTER_LOOP_C_93 : begin
        fsm_output = 8'b01100001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_94;
      end
      LOAD_DATA_OUTER_LOOP_C_94 : begin
        fsm_output = 8'b01100010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_95;
      end
      LOAD_DATA_OUTER_LOOP_C_95 : begin
        fsm_output = 8'b01100011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_96;
      end
      LOAD_DATA_OUTER_LOOP_C_96 : begin
        fsm_output = 8'b01100100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_97;
      end
      LOAD_DATA_OUTER_LOOP_C_97 : begin
        fsm_output = 8'b01100101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_98;
      end
      LOAD_DATA_OUTER_LOOP_C_98 : begin
        fsm_output = 8'b01100110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_99;
      end
      LOAD_DATA_OUTER_LOOP_C_99 : begin
        fsm_output = 8'b01100111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_100;
      end
      LOAD_DATA_OUTER_LOOP_C_100 : begin
        fsm_output = 8'b01101000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_101;
      end
      LOAD_DATA_OUTER_LOOP_C_101 : begin
        fsm_output = 8'b01101001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_102;
      end
      LOAD_DATA_OUTER_LOOP_C_102 : begin
        fsm_output = 8'b01101010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_103;
      end
      LOAD_DATA_OUTER_LOOP_C_103 : begin
        fsm_output = 8'b01101011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_104;
      end
      LOAD_DATA_OUTER_LOOP_C_104 : begin
        fsm_output = 8'b01101100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_105;
      end
      LOAD_DATA_OUTER_LOOP_C_105 : begin
        fsm_output = 8'b01101101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_106;
      end
      LOAD_DATA_OUTER_LOOP_C_106 : begin
        fsm_output = 8'b01101110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_107;
      end
      LOAD_DATA_OUTER_LOOP_C_107 : begin
        fsm_output = 8'b01101111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_108;
      end
      LOAD_DATA_OUTER_LOOP_C_108 : begin
        fsm_output = 8'b01110000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_109;
      end
      LOAD_DATA_OUTER_LOOP_C_109 : begin
        fsm_output = 8'b01110001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_110;
      end
      LOAD_DATA_OUTER_LOOP_C_110 : begin
        fsm_output = 8'b01110010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_111;
      end
      LOAD_DATA_OUTER_LOOP_C_111 : begin
        fsm_output = 8'b01110011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_112;
      end
      LOAD_DATA_OUTER_LOOP_C_112 : begin
        fsm_output = 8'b01110100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_113;
      end
      LOAD_DATA_OUTER_LOOP_C_113 : begin
        fsm_output = 8'b01110101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_114;
      end
      LOAD_DATA_OUTER_LOOP_C_114 : begin
        fsm_output = 8'b01110110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_115;
      end
      LOAD_DATA_OUTER_LOOP_C_115 : begin
        fsm_output = 8'b01110111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_116;
      end
      LOAD_DATA_OUTER_LOOP_C_116 : begin
        fsm_output = 8'b01111000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_117;
      end
      LOAD_DATA_OUTER_LOOP_C_117 : begin
        fsm_output = 8'b01111001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_118;
      end
      LOAD_DATA_OUTER_LOOP_C_118 : begin
        fsm_output = 8'b01111010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_119;
      end
      LOAD_DATA_OUTER_LOOP_C_119 : begin
        fsm_output = 8'b01111011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_120;
      end
      LOAD_DATA_OUTER_LOOP_C_120 : begin
        fsm_output = 8'b01111100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_121;
      end
      LOAD_DATA_OUTER_LOOP_C_121 : begin
        fsm_output = 8'b01111101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_122;
      end
      LOAD_DATA_OUTER_LOOP_C_122 : begin
        fsm_output = 8'b01111110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_123;
      end
      LOAD_DATA_OUTER_LOOP_C_123 : begin
        fsm_output = 8'b01111111;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_124;
      end
      LOAD_DATA_OUTER_LOOP_C_124 : begin
        fsm_output = 8'b10000000;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_125;
      end
      LOAD_DATA_OUTER_LOOP_C_125 : begin
        fsm_output = 8'b10000001;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_126;
      end
      LOAD_DATA_OUTER_LOOP_C_126 : begin
        fsm_output = 8'b10000010;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_127;
      end
      LOAD_DATA_OUTER_LOOP_C_127 : begin
        fsm_output = 8'b10000011;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_128;
      end
      LOAD_DATA_OUTER_LOOP_C_128 : begin
        fsm_output = 8'b10000100;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_129;
      end
      LOAD_DATA_OUTER_LOOP_C_129 : begin
        fsm_output = 8'b10000101;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_130;
      end
      LOAD_DATA_OUTER_LOOP_C_130 : begin
        fsm_output = 8'b10000110;
        state_var_NS = LOAD_DATA_OUTER_LOOP_C_131;
      end
      LOAD_DATA_OUTER_LOOP_C_131 : begin
        fsm_output = 8'b10000111;
        if ( LOAD_DATA_OUTER_LOOP_C_131_tr0 ) begin
          state_var_NS = LOAD_BATCH_LOOP_C_1;
        end
        else begin
          state_var_NS = LOAD_DATA_OUTER_LOOP_C_0;
        end
      end
      LOAD_BATCH_LOOP_C_1 : begin
        fsm_output = 8'b10001000;
        if ( LOAD_BATCH_LOOP_C_1_tr0 ) begin
          state_var_NS = LOAD_BATCH_LOOP_C_0;
        end
        else begin
          state_var_NS = PROCESS_DONE_LOOP_C_0;
        end
      end
      PROCESS_DONE_LOOP_C_0 : begin
        fsm_output = 8'b10001001;
        state_var_NS = PROCESS_DONE_LOOP_C_0;
      end
      // WAIT_FOR_CONFIG_LOOP_C_0
      default : begin
        fsm_output = 8'b00000000;
        if ( WAIT_FOR_CONFIG_LOOP_C_0_tr0 ) begin
          state_var_NS = WAIT_FOR_CONFIG_LOOP_C_0;
        end
        else begin
          state_var_NS = load_input_rlp_C_0;
        end
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= WAIT_FOR_CONFIG_LOOP_C_0;
    end
    else if ( load_input_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_staller
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_staller (
  load_input_wen, dma_read_ctrl_Push_mioi_wen_comp, dma_read_chnl_Pop_mioi_wen_comp,
      input_ready_channel_Pop_mioi_wen_comp, plm_in_cnsi_wen_comp
);
  output load_input_wen;
  input dma_read_ctrl_Push_mioi_wen_comp;
  input dma_read_chnl_Pop_mioi_wen_comp;
  input input_ready_channel_Pop_mioi_wen_comp;
  input plm_in_cnsi_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign load_input_wen = dma_read_ctrl_Push_mioi_wen_comp & dma_read_chnl_Pop_mioi_wen_comp
      & input_ready_channel_Pop_mioi_wen_comp & plm_in_cnsi_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi_plm_in_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi_plm_in_wait_dp (
  clk, rst, plm_in_cnsi_oswt, plm_in_cnsi_wen_comp, plm_in_cnsi_biwt, plm_in_cnsi_bdwt,
      plm_in_cnsi_bcwt
);
  input clk;
  input rst;
  input plm_in_cnsi_oswt;
  output plm_in_cnsi_wen_comp;
  input plm_in_cnsi_biwt;
  input plm_in_cnsi_bdwt;
  output plm_in_cnsi_bcwt;
  reg plm_in_cnsi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cnsi_wen_comp = (~ plm_in_cnsi_oswt) | plm_in_cnsi_biwt | plm_in_cnsi_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      plm_in_cnsi_bcwt <= 1'b0;
    end
    else begin
      plm_in_cnsi_bcwt <= ~((~(plm_in_cnsi_bcwt | plm_in_cnsi_biwt)) | plm_in_cnsi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi_plm_in_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi_plm_in_wait_ctrl
    (
  load_input_wen, plm_in_cnsi_oswt, plm_in_cnsi_irdy, plm_in_cnsi_biwt, plm_in_cnsi_bdwt,
      plm_in_cnsi_bcwt, plm_in_cnsi_ivld_load_input_sct
);
  input load_input_wen;
  input plm_in_cnsi_oswt;
  input plm_in_cnsi_irdy;
  output plm_in_cnsi_biwt;
  output plm_in_cnsi_bdwt;
  input plm_in_cnsi_bcwt;
  output plm_in_cnsi_ivld_load_input_sct;


  // Interconnect Declarations
  wire plm_in_cnsi_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign plm_in_cnsi_bdwt = plm_in_cnsi_oswt & load_input_wen;
  assign plm_in_cnsi_biwt = plm_in_cnsi_ogwt & plm_in_cnsi_irdy;
  assign plm_in_cnsi_ogwt = plm_in_cnsi_oswt & (~ plm_in_cnsi_bcwt);
  assign plm_in_cnsi_ivld_load_input_sct = plm_in_cnsi_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_input_ready_channel_Pop_mioi_input_ready_channel_Pop_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_input_ready_channel_Pop_mioi_input_ready_channel_Pop_mio_wait_dp
    (
  clk, rst, input_ready_channel_Pop_mioi_oswt, input_ready_channel_Pop_mioi_wen_comp,
      input_ready_channel_Pop_mioi_biwt, input_ready_channel_Pop_mioi_bdwt, input_ready_channel_Pop_mioi_bcwt
);
  input clk;
  input rst;
  input input_ready_channel_Pop_mioi_oswt;
  output input_ready_channel_Pop_mioi_wen_comp;
  input input_ready_channel_Pop_mioi_biwt;
  input input_ready_channel_Pop_mioi_bdwt;
  output input_ready_channel_Pop_mioi_bcwt;
  reg input_ready_channel_Pop_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign input_ready_channel_Pop_mioi_wen_comp = (~ input_ready_channel_Pop_mioi_oswt)
      | input_ready_channel_Pop_mioi_biwt | input_ready_channel_Pop_mioi_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      input_ready_channel_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      input_ready_channel_Pop_mioi_bcwt <= ~((~(input_ready_channel_Pop_mioi_bcwt
          | input_ready_channel_Pop_mioi_biwt)) | input_ready_channel_Pop_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_input_ready_channel_Pop_mioi_input_ready_channel_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_input_ready_channel_Pop_mioi_input_ready_channel_Pop_mio_wait_ctrl
    (
  load_input_wen, input_ready_channel_Pop_mioi_oswt, input_ready_channel_Pop_mioi_biwt,
      input_ready_channel_Pop_mioi_bdwt, input_ready_channel_Pop_mioi_bcwt, input_ready_channel_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct,
      input_ready_channel_Pop_mioi_ccs_ccore_done_sync_vld, input_ready_channel_Pop_mioi_oswt_pff
);
  input load_input_wen;
  input input_ready_channel_Pop_mioi_oswt;
  output input_ready_channel_Pop_mioi_biwt;
  output input_ready_channel_Pop_mioi_bdwt;
  input input_ready_channel_Pop_mioi_bcwt;
  output input_ready_channel_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct;
  input input_ready_channel_Pop_mioi_ccs_ccore_done_sync_vld;
  input input_ready_channel_Pop_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign input_ready_channel_Pop_mioi_bdwt = input_ready_channel_Pop_mioi_oswt &
      load_input_wen;
  assign input_ready_channel_Pop_mioi_biwt = input_ready_channel_Pop_mioi_oswt &
      (~ input_ready_channel_Pop_mioi_bcwt) & input_ready_channel_Pop_mioi_ccs_ccore_done_sync_vld;
  assign input_ready_channel_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct = input_ready_channel_Pop_mioi_oswt_pff
      & load_input_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp
    (
  clk, rst, dma_read_chnl_Pop_mioi_oswt, dma_read_chnl_Pop_mioi_wen_comp, dma_read_chnl_Pop_mioi_return_rsc_z_mxwt,
      dma_read_chnl_Pop_mioi_return_rsc_z, dma_read_chnl_Pop_mioi_biwt, dma_read_chnl_Pop_mioi_bdwt,
      dma_read_chnl_Pop_mioi_bcwt
);
  input clk;
  input rst;
  input dma_read_chnl_Pop_mioi_oswt;
  output dma_read_chnl_Pop_mioi_wen_comp;
  output [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt;
  input [63:0] dma_read_chnl_Pop_mioi_return_rsc_z;
  input dma_read_chnl_Pop_mioi_biwt;
  input dma_read_chnl_Pop_mioi_bdwt;
  output dma_read_chnl_Pop_mioi_bcwt;
  reg dma_read_chnl_Pop_mioi_bcwt;


  // Interconnect Declarations
  reg [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_bfwt_31_0;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_chnl_Pop_mioi_wen_comp = (~ dma_read_chnl_Pop_mioi_oswt) | dma_read_chnl_Pop_mioi_biwt
      | dma_read_chnl_Pop_mioi_bcwt;
  assign dma_read_chnl_Pop_mioi_return_rsc_z_mxwt = MUX_v_32_2_2((dma_read_chnl_Pop_mioi_return_rsc_z[31:0]),
      dma_read_chnl_Pop_mioi_return_rsc_z_bfwt_31_0, dma_read_chnl_Pop_mioi_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_chnl_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_read_chnl_Pop_mioi_bcwt <= ~((~(dma_read_chnl_Pop_mioi_bcwt | dma_read_chnl_Pop_mioi_biwt))
          | dma_read_chnl_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( dma_read_chnl_Pop_mioi_biwt ) begin
      dma_read_chnl_Pop_mioi_return_rsc_z_bfwt_31_0 <= dma_read_chnl_Pop_mioi_return_rsc_z[31:0];
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl
    (
  load_input_wen, dma_read_chnl_Pop_mioi_oswt, dma_read_chnl_Pop_mioi_biwt, dma_read_chnl_Pop_mioi_bdwt,
      dma_read_chnl_Pop_mioi_bcwt, dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct,
      dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld, dma_read_chnl_Pop_mioi_oswt_pff
);
  input load_input_wen;
  input dma_read_chnl_Pop_mioi_oswt;
  output dma_read_chnl_Pop_mioi_biwt;
  output dma_read_chnl_Pop_mioi_bdwt;
  input dma_read_chnl_Pop_mioi_bcwt;
  output dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct;
  input dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld;
  input dma_read_chnl_Pop_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dma_read_chnl_Pop_mioi_bdwt = dma_read_chnl_Pop_mioi_oswt & load_input_wen;
  assign dma_read_chnl_Pop_mioi_biwt = dma_read_chnl_Pop_mioi_oswt & (~ dma_read_chnl_Pop_mioi_bcwt)
      & dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld;
  assign dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct = dma_read_chnl_Pop_mioi_oswt_pff
      & load_input_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp
    (
  clk, rst, dma_read_ctrl_Push_mioi_oswt, dma_read_ctrl_Push_mioi_wen_comp, dma_read_ctrl_Push_mioi_biwt,
      dma_read_ctrl_Push_mioi_bdwt, dma_read_ctrl_Push_mioi_bcwt
);
  input clk;
  input rst;
  input dma_read_ctrl_Push_mioi_oswt;
  output dma_read_ctrl_Push_mioi_wen_comp;
  input dma_read_ctrl_Push_mioi_biwt;
  input dma_read_ctrl_Push_mioi_bdwt;
  output dma_read_ctrl_Push_mioi_bcwt;
  reg dma_read_ctrl_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign dma_read_ctrl_Push_mioi_wen_comp = (~ dma_read_ctrl_Push_mioi_oswt) | dma_read_ctrl_Push_mioi_biwt
      | dma_read_ctrl_Push_mioi_bcwt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_read_ctrl_Push_mioi_bcwt <= ~((~(dma_read_ctrl_Push_mioi_bcwt | dma_read_ctrl_Push_mioi_biwt))
          | dma_read_ctrl_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl
    (
  load_input_wen, dma_read_ctrl_Push_mioi_oswt, dma_read_ctrl_Push_mioi_biwt, dma_read_ctrl_Push_mioi_bdwt,
      dma_read_ctrl_Push_mioi_bcwt, dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_input_sct,
      dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld, dma_read_ctrl_Push_mioi_oswt_pff
);
  input load_input_wen;
  input dma_read_ctrl_Push_mioi_oswt;
  output dma_read_ctrl_Push_mioi_biwt;
  output dma_read_ctrl_Push_mioi_bdwt;
  input dma_read_ctrl_Push_mioi_bcwt;
  output dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_input_sct;
  input dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  input dma_read_ctrl_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign dma_read_ctrl_Push_mioi_bdwt = dma_read_ctrl_Push_mioi_oswt & load_input_wen;
  assign dma_read_ctrl_Push_mioi_biwt = dma_read_ctrl_Push_mioi_oswt & (~ dma_read_ctrl_Push_mioi_bcwt)
      & dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  assign dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_input_sct = dma_read_ctrl_Push_mioi_oswt_pff
      & load_input_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_config_accelerator_config_accelerator_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_config_accelerator_config_accelerator_fsm (
  clk, rst, fsm_output, CONFIG_LOOP_C_0_tr0
);
  input clk;
  input rst;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;
  input CONFIG_LOOP_C_0_tr0;


  // FSM State Type Declaration for esp_acc_softmax_softmax_config_accelerator_config_accelerator_fsm_1
  parameter
    config_accelerator_rlp_C_0 = 2'd0,
    CONFIG_LOOP_C_0 = 2'd1,
    CONFIG_DONE_LOOP_C_0 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_softmax_softmax_config_accelerator_config_accelerator_fsm_1
    case (state_var)
      CONFIG_LOOP_C_0 : begin
        fsm_output = 3'b010;
        if ( CONFIG_LOOP_C_0_tr0 ) begin
          state_var_NS = CONFIG_LOOP_C_0;
        end
        else begin
          state_var_NS = CONFIG_DONE_LOOP_C_0;
        end
      end
      CONFIG_DONE_LOOP_C_0 : begin
        fsm_output = 3'b100;
        state_var_NS = CONFIG_DONE_LOOP_C_0;
      end
      // config_accelerator_rlp_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = CONFIG_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= config_accelerator_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi (
  clk, rst, plm_out_cns_dat, plm_out_cns_vld, plm_out_cns_rdy, store_output_wen,
      plm_out_cnsi_oswt, plm_out_cnsi_wen_comp, plm_out_cnsi_idat_mxwt
);
  input clk;
  input rst;
  input [4095:0] plm_out_cns_dat;
  input plm_out_cns_vld;
  output plm_out_cns_rdy;
  input store_output_wen;
  input plm_out_cnsi_oswt;
  output plm_out_cnsi_wen_comp;
  output [4095:0] plm_out_cnsi_idat_mxwt;


  // Interconnect Declarations
  wire plm_out_cnsi_biwt;
  wire plm_out_cnsi_bdwt;
  wire plm_out_cnsi_bcwt;
  wire plm_out_cnsi_irdy_store_output_sct;
  wire plm_out_cnsi_ivld;
  wire [4095:0] plm_out_cnsi_idat;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_ccs_in_wait_v1 #(.rscid(32'sd42),
  .width(32'sd4096)) plm_out_cnsi (
      .rdy(plm_out_cns_rdy),
      .vld(plm_out_cns_vld),
      .dat(plm_out_cns_dat),
      .irdy(plm_out_cnsi_irdy_store_output_sct),
      .ivld(plm_out_cnsi_ivld),
      .idat(plm_out_cnsi_idat)
    );
  esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_plm_out_wait_ctrl
      softmax_store_output_store_output_plm_out_cnsi_plm_out_wait_ctrl_inst (
      .store_output_wen(store_output_wen),
      .plm_out_cnsi_oswt(plm_out_cnsi_oswt),
      .plm_out_cnsi_biwt(plm_out_cnsi_biwt),
      .plm_out_cnsi_bdwt(plm_out_cnsi_bdwt),
      .plm_out_cnsi_bcwt(plm_out_cnsi_bcwt),
      .plm_out_cnsi_irdy_store_output_sct(plm_out_cnsi_irdy_store_output_sct),
      .plm_out_cnsi_ivld(plm_out_cnsi_ivld)
    );
  esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi_plm_out_wait_dp
      softmax_store_output_store_output_plm_out_cnsi_plm_out_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_out_cnsi_oswt(plm_out_cnsi_oswt),
      .plm_out_cnsi_wen_comp(plm_out_cnsi_wen_comp),
      .plm_out_cnsi_idat_mxwt(plm_out_cnsi_idat_mxwt),
      .plm_out_cnsi_biwt(plm_out_cnsi_biwt),
      .plm_out_cnsi_bdwt(plm_out_cnsi_bdwt),
      .plm_out_cnsi_bcwt(plm_out_cnsi_bcwt),
      .plm_out_cnsi_idat(plm_out_cnsi_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi
    (
  clk, rst, dma_write_chnl_val, dma_write_chnl_rdy, dma_write_chnl_msg, store_output_wen,
      dma_write_chnl_Push_mioi_oswt, dma_write_chnl_Push_mioi_wen_comp, dma_write_chnl_Push_mioi_m_rsc_dat_store_output,
      dma_write_chnl_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;
  input store_output_wen;
  input dma_write_chnl_Push_mioi_oswt;
  output dma_write_chnl_Push_mioi_wen_comp;
  input [63:0] dma_write_chnl_Push_mioi_m_rsc_dat_store_output;
  input dma_write_chnl_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire [63:0] dma_write_chnl_Push_mioi_m_rsc_dat;
  wire dma_write_chnl_Push_mioi_biwt;
  wire dma_write_chnl_Push_mioi_bdwt;
  wire dma_write_chnl_Push_mioi_bcwt;
  wire dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld;
  wire dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [63:0] nl_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp_inst_dma_write_chnl_Push_mioi_m_rsc_dat_store_output;
  assign nl_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp_inst_dma_write_chnl_Push_mioi_m_rsc_dat_store_output
      = {32'b11011110101011011011111011101111 , (dma_write_chnl_Push_mioi_m_rsc_dat_store_output[31:0])};
  esp_acc_softmax_Connections_OutBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Push
      dma_write_chnl_Push_mioi (
      .this_val(dma_write_chnl_val),
      .this_rdy(dma_write_chnl_rdy),
      .this_msg(dma_write_chnl_msg),
      .m_rsc_dat(dma_write_chnl_Push_mioi_m_rsc_dat),
      .ccs_ccore_start_rsc_dat(dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_iff),
      .ccs_ccore_done_sync_vld(dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl
      softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl_inst
      (
      .store_output_wen(store_output_wen),
      .dma_write_chnl_Push_mioi_oswt(dma_write_chnl_Push_mioi_oswt),
      .dma_write_chnl_Push_mioi_biwt(dma_write_chnl_Push_mioi_biwt),
      .dma_write_chnl_Push_mioi_bdwt(dma_write_chnl_Push_mioi_bdwt),
      .dma_write_chnl_Push_mioi_bcwt(dma_write_chnl_Push_mioi_bcwt),
      .dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld(dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld),
      .dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff(dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_iff),
      .dma_write_chnl_Push_mioi_oswt_pff(dma_write_chnl_Push_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp
      softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_chnl_Push_mioi_oswt(dma_write_chnl_Push_mioi_oswt),
      .dma_write_chnl_Push_mioi_wen_comp(dma_write_chnl_Push_mioi_wen_comp),
      .dma_write_chnl_Push_mioi_m_rsc_dat_store_output(nl_softmax_store_output_store_output_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp_inst_dma_write_chnl_Push_mioi_m_rsc_dat_store_output[63:0]),
      .dma_write_chnl_Push_mioi_m_rsc_dat(dma_write_chnl_Push_mioi_m_rsc_dat),
      .dma_write_chnl_Push_mioi_biwt(dma_write_chnl_Push_mioi_biwt),
      .dma_write_chnl_Push_mioi_bdwt(dma_write_chnl_Push_mioi_bdwt),
      .dma_write_chnl_Push_mioi_bcwt(dma_write_chnl_Push_mioi_bcwt),
      .dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_pff(dma_write_chnl_Push_mioi_m_rsc_dat_store_output_sct_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi
    (
  clk, rst, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg, store_output_wen,
      dma_write_ctrl_Push_mioi_oswt, dma_write_ctrl_Push_mioi_wen_comp, dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output,
      dma_write_ctrl_Push_mioi_m_length_rsc_dat_store_output, dma_write_ctrl_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  input store_output_wen;
  input dma_write_ctrl_Push_mioi_oswt;
  output dma_write_ctrl_Push_mioi_wen_comp;
  input [31:0] dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output;
  input [31:0] dma_write_ctrl_Push_mioi_m_length_rsc_dat_store_output;
  input dma_write_ctrl_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire dma_write_ctrl_Push_mioi_biwt;
  wire dma_write_ctrl_Push_mioi_bdwt;
  wire dma_write_ctrl_Push_mioi_bcwt;
  wire dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_output_sct;
  wire dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push  dma_write_ctrl_Push_mioi
      (
      .this_val(dma_write_ctrl_val),
      .this_rdy(dma_write_ctrl_rdy),
      .this_msg(dma_write_ctrl_msg),
      .m_index_rsc_dat(dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output),
      .m_length_rsc_dat(dma_write_ctrl_Push_mioi_m_length_rsc_dat_store_output),
      .ccs_ccore_start_rsc_dat(dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_output_sct),
      .ccs_ccore_done_sync_vld(dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl
      softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl_inst
      (
      .store_output_wen(store_output_wen),
      .dma_write_ctrl_Push_mioi_oswt(dma_write_ctrl_Push_mioi_oswt),
      .dma_write_ctrl_Push_mioi_biwt(dma_write_ctrl_Push_mioi_biwt),
      .dma_write_ctrl_Push_mioi_bdwt(dma_write_ctrl_Push_mioi_bdwt),
      .dma_write_ctrl_Push_mioi_bcwt(dma_write_ctrl_Push_mioi_bcwt),
      .dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_output_sct(dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_store_output_sct),
      .dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld(dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .dma_write_ctrl_Push_mioi_oswt_pff(dma_write_ctrl_Push_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp
      softmax_store_output_store_output_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_ctrl_Push_mioi_oswt(dma_write_ctrl_Push_mioi_oswt),
      .dma_write_ctrl_Push_mioi_wen_comp(dma_write_ctrl_Push_mioi_wen_comp),
      .dma_write_ctrl_Push_mioi_biwt(dma_write_ctrl_Push_mioi_biwt),
      .dma_write_ctrl_Push_mioi_bdwt(dma_write_ctrl_Push_mioi_bdwt),
      .dma_write_ctrl_Push_mioi_bcwt(dma_write_ctrl_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output_output_ready_channel_Push_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output_output_ready_channel_Push_mioi
    (
  clk, rst, output_ready_channel_val, output_ready_channel_rdy, output_ready_channel_msg,
      store_output_wen, output_ready_channel_Push_mioi_oswt, output_ready_channel_Push_mioi_wen_comp,
      output_ready_channel_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output output_ready_channel_val;
  input output_ready_channel_rdy;
  output output_ready_channel_msg;
  input store_output_wen;
  input output_ready_channel_Push_mioi_oswt;
  output output_ready_channel_Push_mioi_wen_comp;
  input output_ready_channel_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire output_ready_channel_Push_mioi_biwt;
  wire output_ready_channel_Push_mioi_bdwt;
  wire output_ready_channel_Push_mioi_bcwt;
  wire output_ready_channel_Push_mioi_ccs_ccore_start_rsc_dat_store_output_sct;
  wire output_ready_channel_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_Connections_Combinational_bool_Connections_SYN_PORT_Push  output_ready_channel_Push_mioi
      (
      .this_val(output_ready_channel_val),
      .this_rdy(output_ready_channel_rdy),
      .this_msg(output_ready_channel_msg),
      .ccs_ccore_start_rsc_dat(output_ready_channel_Push_mioi_ccs_ccore_start_rsc_dat_store_output_sct),
      .ccs_ccore_done_sync_vld(output_ready_channel_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_store_output_store_output_output_ready_channel_Push_mioi_output_ready_channel_Push_mio_wait_ctrl
      softmax_store_output_store_output_output_ready_channel_Push_mioi_output_ready_channel_Push_mio_wait_ctrl_inst
      (
      .store_output_wen(store_output_wen),
      .output_ready_channel_Push_mioi_oswt(output_ready_channel_Push_mioi_oswt),
      .output_ready_channel_Push_mioi_biwt(output_ready_channel_Push_mioi_biwt),
      .output_ready_channel_Push_mioi_bdwt(output_ready_channel_Push_mioi_bdwt),
      .output_ready_channel_Push_mioi_bcwt(output_ready_channel_Push_mioi_bcwt),
      .output_ready_channel_Push_mioi_ccs_ccore_start_rsc_dat_store_output_sct(output_ready_channel_Push_mioi_ccs_ccore_start_rsc_dat_store_output_sct),
      .output_ready_channel_Push_mioi_ccs_ccore_done_sync_vld(output_ready_channel_Push_mioi_ccs_ccore_done_sync_vld),
      .output_ready_channel_Push_mioi_oswt_pff(output_ready_channel_Push_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_store_output_store_output_output_ready_channel_Push_mioi_output_ready_channel_Push_mio_wait_dp
      softmax_store_output_store_output_output_ready_channel_Push_mioi_output_ready_channel_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .output_ready_channel_Push_mioi_oswt(output_ready_channel_Push_mioi_oswt),
      .output_ready_channel_Push_mioi_wen_comp(output_ready_channel_Push_mioi_wen_comp),
      .output_ready_channel_Push_mioi_biwt(output_ready_channel_Push_mioi_biwt),
      .output_ready_channel_Push_mioi_bdwt(output_ready_channel_Push_mioi_bdwt),
      .output_ready_channel_Push_mioi_bcwt(output_ready_channel_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi (
  clk, rst, plm_out_cns_dat, plm_out_cns_vld, plm_out_cns_rdy, compute_kernel_wen,
      plm_out_cnsi_oswt, plm_out_cnsi_wen_comp, plm_out_cnsi_idat
);
  input clk;
  input rst;
  output [4095:0] plm_out_cns_dat;
  output plm_out_cns_vld;
  input plm_out_cns_rdy;
  input compute_kernel_wen;
  input plm_out_cnsi_oswt;
  output plm_out_cnsi_wen_comp;
  input [4095:0] plm_out_cnsi_idat;


  // Interconnect Declarations
  wire plm_out_cnsi_irdy;
  wire plm_out_cnsi_biwt;
  wire plm_out_cnsi_bdwt;
  wire plm_out_cnsi_bcwt;
  wire plm_out_cnsi_ivld_compute_kernel_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_ccs_out_wait_v1 #(.rscid(32'sd37),
  .width(32'sd4096)) plm_out_cnsi (
      .irdy(plm_out_cnsi_irdy),
      .ivld(plm_out_cnsi_ivld_compute_kernel_sct),
      .idat(plm_out_cnsi_idat),
      .rdy(plm_out_cns_rdy),
      .vld(plm_out_cns_vld),
      .dat(plm_out_cns_dat)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi_plm_out_wait_ctrl
      softmax_compute_kernel_compute_kernel_plm_out_cnsi_plm_out_wait_ctrl_inst (
      .compute_kernel_wen(compute_kernel_wen),
      .plm_out_cnsi_oswt(plm_out_cnsi_oswt),
      .plm_out_cnsi_irdy(plm_out_cnsi_irdy),
      .plm_out_cnsi_biwt(plm_out_cnsi_biwt),
      .plm_out_cnsi_bdwt(plm_out_cnsi_bdwt),
      .plm_out_cnsi_bcwt(plm_out_cnsi_bcwt),
      .plm_out_cnsi_ivld_compute_kernel_sct(plm_out_cnsi_ivld_compute_kernel_sct)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi_plm_out_wait_dp
      softmax_compute_kernel_compute_kernel_plm_out_cnsi_plm_out_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_out_cnsi_oswt(plm_out_cnsi_oswt),
      .plm_out_cnsi_wen_comp(plm_out_cnsi_wen_comp),
      .plm_out_cnsi_biwt(plm_out_cnsi_biwt),
      .plm_out_cnsi_bdwt(plm_out_cnsi_bdwt),
      .plm_out_cnsi_bcwt(plm_out_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi (
  clk, rst, plm_in_cns_dat, plm_in_cns_vld, plm_in_cns_rdy, compute_kernel_wen, plm_in_cnsi_oswt,
      plm_in_cnsi_wen_comp, plm_in_cnsi_idat_mxwt
);
  input clk;
  input rst;
  input [4095:0] plm_in_cns_dat;
  input plm_in_cns_vld;
  output plm_in_cns_rdy;
  input compute_kernel_wen;
  input plm_in_cnsi_oswt;
  output plm_in_cnsi_wen_comp;
  output [4095:0] plm_in_cnsi_idat_mxwt;


  // Interconnect Declarations
  wire plm_in_cnsi_biwt;
  wire plm_in_cnsi_bdwt;
  wire plm_in_cnsi_bcwt;
  wire plm_in_cnsi_irdy_compute_kernel_sct;
  wire plm_in_cnsi_ivld;
  wire [4095:0] plm_in_cnsi_idat;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_ccs_in_wait_v1 #(.rscid(32'sd36),
  .width(32'sd4096)) plm_in_cnsi (
      .rdy(plm_in_cns_rdy),
      .vld(plm_in_cns_vld),
      .dat(plm_in_cns_dat),
      .irdy(plm_in_cnsi_irdy_compute_kernel_sct),
      .ivld(plm_in_cnsi_ivld),
      .idat(plm_in_cnsi_idat)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_plm_in_wait_ctrl
      softmax_compute_kernel_compute_kernel_plm_in_cnsi_plm_in_wait_ctrl_inst (
      .compute_kernel_wen(compute_kernel_wen),
      .plm_in_cnsi_oswt(plm_in_cnsi_oswt),
      .plm_in_cnsi_biwt(plm_in_cnsi_biwt),
      .plm_in_cnsi_bdwt(plm_in_cnsi_bdwt),
      .plm_in_cnsi_bcwt(plm_in_cnsi_bcwt),
      .plm_in_cnsi_irdy_compute_kernel_sct(plm_in_cnsi_irdy_compute_kernel_sct),
      .plm_in_cnsi_ivld(plm_in_cnsi_ivld)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi_plm_in_wait_dp
      softmax_compute_kernel_compute_kernel_plm_in_cnsi_plm_in_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .plm_in_cnsi_oswt(plm_in_cnsi_oswt),
      .plm_in_cnsi_wen_comp(plm_in_cnsi_wen_comp),
      .plm_in_cnsi_idat_mxwt(plm_in_cnsi_idat_mxwt),
      .plm_in_cnsi_biwt(plm_in_cnsi_biwt),
      .plm_in_cnsi_bdwt(plm_in_cnsi_bdwt),
      .plm_in_cnsi_bcwt(plm_in_cnsi_bcwt),
      .plm_in_cnsi_idat(plm_in_cnsi_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_channel_Pop_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_channel_Pop_mioi
    (
  clk, rst, output_ready_channel_val, output_ready_channel_rdy, output_ready_channel_msg,
      compute_kernel_wen, output_ready_channel_Pop_mioi_oswt, output_ready_channel_Pop_mioi_wen_comp,
      output_ready_channel_Pop_mioi_oswt_pff
);
  input clk;
  input rst;
  input output_ready_channel_val;
  output output_ready_channel_rdy;
  input output_ready_channel_msg;
  input compute_kernel_wen;
  input output_ready_channel_Pop_mioi_oswt;
  output output_ready_channel_Pop_mioi_wen_comp;
  input output_ready_channel_Pop_mioi_oswt_pff;


  // Interconnect Declarations
  wire output_ready_channel_Pop_mioi_return_rsc_z;
  wire output_ready_channel_Pop_mioi_biwt;
  wire output_ready_channel_Pop_mioi_bdwt;
  wire output_ready_channel_Pop_mioi_bcwt;
  wire output_ready_channel_Pop_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct;
  wire output_ready_channel_Pop_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_Connections_Combinational_bool_Connections_SYN_PORT_Pop  output_ready_channel_Pop_mioi
      (
      .this_val(output_ready_channel_val),
      .this_rdy(output_ready_channel_rdy),
      .this_msg(output_ready_channel_msg),
      .return_rsc_z(output_ready_channel_Pop_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(output_ready_channel_Pop_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct),
      .ccs_ccore_done_sync_vld(output_ready_channel_Pop_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_channel_Pop_mioi_output_ready_channel_Pop_mio_wait_ctrl
      softmax_compute_kernel_compute_kernel_output_ready_channel_Pop_mioi_output_ready_channel_Pop_mio_wait_ctrl_inst
      (
      .compute_kernel_wen(compute_kernel_wen),
      .output_ready_channel_Pop_mioi_oswt(output_ready_channel_Pop_mioi_oswt),
      .output_ready_channel_Pop_mioi_biwt(output_ready_channel_Pop_mioi_biwt),
      .output_ready_channel_Pop_mioi_bdwt(output_ready_channel_Pop_mioi_bdwt),
      .output_ready_channel_Pop_mioi_bcwt(output_ready_channel_Pop_mioi_bcwt),
      .output_ready_channel_Pop_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct(output_ready_channel_Pop_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct),
      .output_ready_channel_Pop_mioi_ccs_ccore_done_sync_vld(output_ready_channel_Pop_mioi_ccs_ccore_done_sync_vld),
      .output_ready_channel_Pop_mioi_oswt_pff(output_ready_channel_Pop_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_channel_Pop_mioi_output_ready_channel_Pop_mio_wait_dp
      softmax_compute_kernel_compute_kernel_output_ready_channel_Pop_mioi_output_ready_channel_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .output_ready_channel_Pop_mioi_oswt(output_ready_channel_Pop_mioi_oswt),
      .output_ready_channel_Pop_mioi_wen_comp(output_ready_channel_Pop_mioi_wen_comp),
      .output_ready_channel_Pop_mioi_biwt(output_ready_channel_Pop_mioi_biwt),
      .output_ready_channel_Pop_mioi_bdwt(output_ready_channel_Pop_mioi_bdwt),
      .output_ready_channel_Pop_mioi_bcwt(output_ready_channel_Pop_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_channel_Push_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_channel_Push_mioi
    (
  clk, rst, input_ready_channel_val, input_ready_channel_rdy, input_ready_channel_msg,
      compute_kernel_wen, input_ready_channel_Push_mioi_oswt, input_ready_channel_Push_mioi_wen_comp,
      input_ready_channel_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output input_ready_channel_val;
  input input_ready_channel_rdy;
  output input_ready_channel_msg;
  input compute_kernel_wen;
  input input_ready_channel_Push_mioi_oswt;
  output input_ready_channel_Push_mioi_wen_comp;
  input input_ready_channel_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire input_ready_channel_Push_mioi_biwt;
  wire input_ready_channel_Push_mioi_bdwt;
  wire input_ready_channel_Push_mioi_bcwt;
  wire input_ready_channel_Push_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct;
  wire input_ready_channel_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_Connections_Combinational_bool_Connections_SYN_PORT_Push  input_ready_channel_Push_mioi
      (
      .this_val(input_ready_channel_val),
      .this_rdy(input_ready_channel_rdy),
      .this_msg(input_ready_channel_msg),
      .ccs_ccore_start_rsc_dat(input_ready_channel_Push_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct),
      .ccs_ccore_done_sync_vld(input_ready_channel_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_channel_Push_mioi_input_ready_channel_Push_mio_wait_ctrl
      softmax_compute_kernel_compute_kernel_input_ready_channel_Push_mioi_input_ready_channel_Push_mio_wait_ctrl_inst
      (
      .compute_kernel_wen(compute_kernel_wen),
      .input_ready_channel_Push_mioi_oswt(input_ready_channel_Push_mioi_oswt),
      .input_ready_channel_Push_mioi_biwt(input_ready_channel_Push_mioi_biwt),
      .input_ready_channel_Push_mioi_bdwt(input_ready_channel_Push_mioi_bdwt),
      .input_ready_channel_Push_mioi_bcwt(input_ready_channel_Push_mioi_bcwt),
      .input_ready_channel_Push_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct(input_ready_channel_Push_mioi_ccs_ccore_start_rsc_dat_compute_kernel_sct),
      .input_ready_channel_Push_mioi_ccs_ccore_done_sync_vld(input_ready_channel_Push_mioi_ccs_ccore_done_sync_vld),
      .input_ready_channel_Push_mioi_oswt_pff(input_ready_channel_Push_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_channel_Push_mioi_input_ready_channel_Push_mio_wait_dp
      softmax_compute_kernel_compute_kernel_input_ready_channel_Push_mioi_input_ready_channel_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_ready_channel_Push_mioi_oswt(input_ready_channel_Push_mioi_oswt),
      .input_ready_channel_Push_mioi_wen_comp(input_ready_channel_Push_mioi_wen_comp),
      .input_ready_channel_Push_mioi_biwt(input_ready_channel_Push_mioi_biwt),
      .input_ready_channel_Push_mioi_bdwt(input_ready_channel_Push_mioi_bdwt),
      .input_ready_channel_Push_mioi_bcwt(input_ready_channel_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi (
  clk, rst, plm_in_cns_dat, plm_in_cns_vld, plm_in_cns_rdy, load_input_wen, plm_in_cnsi_oswt,
      plm_in_cnsi_wen_comp, plm_in_cnsi_idat
);
  input clk;
  input rst;
  output [4095:0] plm_in_cns_dat;
  output plm_in_cns_vld;
  input plm_in_cns_rdy;
  input load_input_wen;
  input plm_in_cnsi_oswt;
  output plm_in_cnsi_wen_comp;
  input [4095:0] plm_in_cnsi_idat;


  // Interconnect Declarations
  wire plm_in_cnsi_irdy;
  wire plm_in_cnsi_biwt;
  wire plm_in_cnsi_bdwt;
  wire plm_in_cnsi_bcwt;
  wire plm_in_cnsi_ivld_load_input_sct;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_ccs_out_wait_v1 #(.rscid(32'sd35),
  .width(32'sd4096)) plm_in_cnsi (
      .irdy(plm_in_cnsi_irdy),
      .ivld(plm_in_cnsi_ivld_load_input_sct),
      .idat(plm_in_cnsi_idat),
      .rdy(plm_in_cns_rdy),
      .vld(plm_in_cns_vld),
      .dat(plm_in_cns_dat)
    );
  esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi_plm_in_wait_ctrl softmax_load_input_load_input_plm_in_cnsi_plm_in_wait_ctrl_inst
      (
      .load_input_wen(load_input_wen),
      .plm_in_cnsi_oswt(plm_in_cnsi_oswt),
      .plm_in_cnsi_irdy(plm_in_cnsi_irdy),
      .plm_in_cnsi_biwt(plm_in_cnsi_biwt),
      .plm_in_cnsi_bdwt(plm_in_cnsi_bdwt),
      .plm_in_cnsi_bcwt(plm_in_cnsi_bcwt),
      .plm_in_cnsi_ivld_load_input_sct(plm_in_cnsi_ivld_load_input_sct)
    );
  esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi_plm_in_wait_dp softmax_load_input_load_input_plm_in_cnsi_plm_in_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cnsi_oswt(plm_in_cnsi_oswt),
      .plm_in_cnsi_wen_comp(plm_in_cnsi_wen_comp),
      .plm_in_cnsi_biwt(plm_in_cnsi_biwt),
      .plm_in_cnsi_bdwt(plm_in_cnsi_bdwt),
      .plm_in_cnsi_bcwt(plm_in_cnsi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_input_ready_channel_Pop_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_input_ready_channel_Pop_mioi
    (
  clk, rst, input_ready_channel_val, input_ready_channel_rdy, input_ready_channel_msg,
      load_input_wen, input_ready_channel_Pop_mioi_oswt, input_ready_channel_Pop_mioi_wen_comp,
      input_ready_channel_Pop_mioi_oswt_pff
);
  input clk;
  input rst;
  input input_ready_channel_val;
  output input_ready_channel_rdy;
  input input_ready_channel_msg;
  input load_input_wen;
  input input_ready_channel_Pop_mioi_oswt;
  output input_ready_channel_Pop_mioi_wen_comp;
  input input_ready_channel_Pop_mioi_oswt_pff;


  // Interconnect Declarations
  wire input_ready_channel_Pop_mioi_return_rsc_z;
  wire input_ready_channel_Pop_mioi_biwt;
  wire input_ready_channel_Pop_mioi_bdwt;
  wire input_ready_channel_Pop_mioi_bcwt;
  wire input_ready_channel_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct;
  wire input_ready_channel_Pop_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_Connections_Combinational_bool_Connections_SYN_PORT_Pop  input_ready_channel_Pop_mioi
      (
      .this_val(input_ready_channel_val),
      .this_rdy(input_ready_channel_rdy),
      .this_msg(input_ready_channel_msg),
      .return_rsc_z(input_ready_channel_Pop_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(input_ready_channel_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct),
      .ccs_ccore_done_sync_vld(input_ready_channel_Pop_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_load_input_load_input_input_ready_channel_Pop_mioi_input_ready_channel_Pop_mio_wait_ctrl
      softmax_load_input_load_input_input_ready_channel_Pop_mioi_input_ready_channel_Pop_mio_wait_ctrl_inst
      (
      .load_input_wen(load_input_wen),
      .input_ready_channel_Pop_mioi_oswt(input_ready_channel_Pop_mioi_oswt),
      .input_ready_channel_Pop_mioi_biwt(input_ready_channel_Pop_mioi_biwt),
      .input_ready_channel_Pop_mioi_bdwt(input_ready_channel_Pop_mioi_bdwt),
      .input_ready_channel_Pop_mioi_bcwt(input_ready_channel_Pop_mioi_bcwt),
      .input_ready_channel_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct(input_ready_channel_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct),
      .input_ready_channel_Pop_mioi_ccs_ccore_done_sync_vld(input_ready_channel_Pop_mioi_ccs_ccore_done_sync_vld),
      .input_ready_channel_Pop_mioi_oswt_pff(input_ready_channel_Pop_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_load_input_load_input_input_ready_channel_Pop_mioi_input_ready_channel_Pop_mio_wait_dp
      softmax_load_input_load_input_input_ready_channel_Pop_mioi_input_ready_channel_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_ready_channel_Pop_mioi_oswt(input_ready_channel_Pop_mioi_oswt),
      .input_ready_channel_Pop_mioi_wen_comp(input_ready_channel_Pop_mioi_wen_comp),
      .input_ready_channel_Pop_mioi_biwt(input_ready_channel_Pop_mioi_biwt),
      .input_ready_channel_Pop_mioi_bdwt(input_ready_channel_Pop_mioi_bdwt),
      .input_ready_channel_Pop_mioi_bcwt(input_ready_channel_Pop_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi (
  clk, rst, dma_read_chnl_val, dma_read_chnl_rdy, dma_read_chnl_msg, load_input_wen,
      dma_read_chnl_Pop_mioi_oswt, dma_read_chnl_Pop_mioi_wen_comp, dma_read_chnl_Pop_mioi_return_rsc_z_mxwt,
      dma_read_chnl_Pop_mioi_oswt_pff
);
  input clk;
  input rst;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  input load_input_wen;
  input dma_read_chnl_Pop_mioi_oswt;
  output dma_read_chnl_Pop_mioi_wen_comp;
  output [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt;
  input dma_read_chnl_Pop_mioi_oswt_pff;


  // Interconnect Declarations
  wire [63:0] dma_read_chnl_Pop_mioi_return_rsc_z;
  wire dma_read_chnl_Pop_mioi_biwt;
  wire dma_read_chnl_Pop_mioi_bdwt;
  wire dma_read_chnl_Pop_mioi_bcwt;
  wire dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct;
  wire dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld;
  wire [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_Connections_InBlocking_sc_dt_sc_bv_64_Connections_SYN_PORT_Pop
      dma_read_chnl_Pop_mioi (
      .this_val(dma_read_chnl_val),
      .this_rdy(dma_read_chnl_rdy),
      .this_msg(dma_read_chnl_msg),
      .return_rsc_z(dma_read_chnl_Pop_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct),
      .ccs_ccore_done_sync_vld(dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl
      softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl_inst
      (
      .load_input_wen(load_input_wen),
      .dma_read_chnl_Pop_mioi_oswt(dma_read_chnl_Pop_mioi_oswt),
      .dma_read_chnl_Pop_mioi_biwt(dma_read_chnl_Pop_mioi_biwt),
      .dma_read_chnl_Pop_mioi_bdwt(dma_read_chnl_Pop_mioi_bdwt),
      .dma_read_chnl_Pop_mioi_bcwt(dma_read_chnl_Pop_mioi_bcwt),
      .dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct(dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_load_input_sct),
      .dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld(dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld),
      .dma_read_chnl_Pop_mioi_oswt_pff(dma_read_chnl_Pop_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp
      softmax_load_input_load_input_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_chnl_Pop_mioi_oswt(dma_read_chnl_Pop_mioi_oswt),
      .dma_read_chnl_Pop_mioi_wen_comp(dma_read_chnl_Pop_mioi_wen_comp),
      .dma_read_chnl_Pop_mioi_return_rsc_z_mxwt(dma_read_chnl_Pop_mioi_return_rsc_z_mxwt_pconst),
      .dma_read_chnl_Pop_mioi_return_rsc_z(dma_read_chnl_Pop_mioi_return_rsc_z),
      .dma_read_chnl_Pop_mioi_biwt(dma_read_chnl_Pop_mioi_biwt),
      .dma_read_chnl_Pop_mioi_bdwt(dma_read_chnl_Pop_mioi_bdwt),
      .dma_read_chnl_Pop_mioi_bcwt(dma_read_chnl_Pop_mioi_bcwt)
    );
  assign dma_read_chnl_Pop_mioi_return_rsc_z_mxwt = dma_read_chnl_Pop_mioi_return_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi (
  clk, rst, dma_read_ctrl_val, dma_read_ctrl_rdy, dma_read_ctrl_msg, load_input_wen,
      dma_read_ctrl_Push_mioi_oswt, dma_read_ctrl_Push_mioi_wen_comp, dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input,
      dma_read_ctrl_Push_mioi_m_length_rsc_dat_load_input, dma_read_ctrl_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  input load_input_wen;
  input dma_read_ctrl_Push_mioi_oswt;
  output dma_read_ctrl_Push_mioi_wen_comp;
  input [31:0] dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input;
  input [31:0] dma_read_ctrl_Push_mioi_m_length_rsc_dat_load_input;
  input dma_read_ctrl_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire dma_read_ctrl_Push_mioi_biwt;
  wire dma_read_ctrl_Push_mioi_bdwt;
  wire dma_read_ctrl_Push_mioi_bcwt;
  wire dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_input_sct;
  wire dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push  dma_read_ctrl_Push_mioi
      (
      .this_val(dma_read_ctrl_val),
      .this_rdy(dma_read_ctrl_rdy),
      .this_msg(dma_read_ctrl_msg),
      .m_index_rsc_dat(dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input),
      .m_length_rsc_dat(dma_read_ctrl_Push_mioi_m_length_rsc_dat_load_input),
      .ccs_ccore_start_rsc_dat(dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_input_sct),
      .ccs_ccore_done_sync_vld(dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl
      softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl_inst
      (
      .load_input_wen(load_input_wen),
      .dma_read_ctrl_Push_mioi_oswt(dma_read_ctrl_Push_mioi_oswt),
      .dma_read_ctrl_Push_mioi_biwt(dma_read_ctrl_Push_mioi_biwt),
      .dma_read_ctrl_Push_mioi_bdwt(dma_read_ctrl_Push_mioi_bdwt),
      .dma_read_ctrl_Push_mioi_bcwt(dma_read_ctrl_Push_mioi_bcwt),
      .dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_input_sct(dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_load_input_sct),
      .dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld(dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .dma_read_ctrl_Push_mioi_oswt_pff(dma_read_ctrl_Push_mioi_oswt_pff)
    );
  esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp
      softmax_load_input_load_input_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_ctrl_Push_mioi_oswt(dma_read_ctrl_Push_mioi_oswt),
      .dma_read_ctrl_Push_mioi_wen_comp(dma_read_ctrl_Push_mioi_wen_comp),
      .dma_read_ctrl_Push_mioi_biwt(dma_read_ctrl_Push_mioi_biwt),
      .dma_read_ctrl_Push_mioi_bdwt(dma_read_ctrl_Push_mioi_bdwt),
      .dma_read_ctrl_Push_mioi_bcwt(dma_read_ctrl_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_config_accelerator
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_config_accelerator (
  clk, rst, conf_done, done
);
  input clk;
  input rst;
  input conf_done;
  output done;
  reg done;


  // Interconnect Declarations
  wire [2:0] fsm_output;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_softmax_config_accelerator_config_accelerator_fsm_inst_CONFIG_LOOP_C_0_tr0;
  assign nl_softmax_config_accelerator_config_accelerator_fsm_inst_CONFIG_LOOP_C_0_tr0
      = ~ conf_done;
  esp_acc_softmax_softmax_config_accelerator_config_accelerator_fsm softmax_config_accelerator_config_accelerator_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .CONFIG_LOOP_C_0_tr0(nl_softmax_config_accelerator_config_accelerator_fsm_inst_CONFIG_LOOP_C_0_tr0[0:0])
    );
  always @(posedge clk) begin
    if ( ~ rst ) begin
      done <= 1'b0;
    end
    else if ( conf_done & (fsm_output[1]) ) begin
      done <= 1'b1;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output_store_output
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output_store_output (
  clk, rst, conf_info, acc_done, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg,
      dma_write_chnl_val, dma_write_chnl_rdy, dma_write_chnl_msg, done, output_ready_channel_val,
      output_ready_channel_rdy, output_ready_channel_msg, plm_out_cns_dat, plm_out_cns_vld,
      plm_out_cns_rdy, STORE_MAIN_LOOP_plm_local_data_rsci_clken_d, STORE_MAIN_LOOP_plm_local_data_rsci_d_d,
      STORE_MAIN_LOOP_plm_local_data_rsci_q_d, STORE_MAIN_LOOP_plm_local_data_rsci_radr_d,
      STORE_MAIN_LOOP_plm_local_data_rsci_wadr_d, STORE_MAIN_LOOP_plm_local_data_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      STORE_MAIN_LOOP_plm_local_data_rsci_we_d_pff
);
  input clk;
  input rst;
  input [63:0] conf_info;
  output acc_done;
  reg acc_done;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;
  input done;
  output output_ready_channel_val;
  input output_ready_channel_rdy;
  output output_ready_channel_msg;
  input [4095:0] plm_out_cns_dat;
  input plm_out_cns_vld;
  output plm_out_cns_rdy;
  output STORE_MAIN_LOOP_plm_local_data_rsci_clken_d;
  output [31:0] STORE_MAIN_LOOP_plm_local_data_rsci_d_d;
  input [31:0] STORE_MAIN_LOOP_plm_local_data_rsci_q_d;
  output [6:0] STORE_MAIN_LOOP_plm_local_data_rsci_radr_d;
  output [6:0] STORE_MAIN_LOOP_plm_local_data_rsci_wadr_d;
  output STORE_MAIN_LOOP_plm_local_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output STORE_MAIN_LOOP_plm_local_data_rsci_we_d_pff;


  // Interconnect Declarations
  wire store_output_wen;
  wire output_ready_channel_Push_mioi_wen_comp;
  wire dma_write_ctrl_Push_mioi_wen_comp;
  wire dma_write_chnl_Push_mioi_wen_comp;
  wire plm_out_cnsi_wen_comp;
  wire [4095:0] plm_out_cnsi_idat_mxwt;
  wire [7:0] fsm_output;
  wire and_dcpl_3;
  wire and_dcpl_5;
  wire and_dcpl_8;
  wire and_dcpl_9;
  wire and_dcpl_10;
  wire and_dcpl_12;
  wire or_dcpl_1;
  wire and_dcpl_14;
  wire and_dcpl_15;
  wire and_dcpl_16;
  wire and_dcpl_17;
  wire and_dcpl_18;
  wire and_dcpl_19;
  wire and_dcpl_20;
  wire and_dcpl_21;
  wire and_dcpl_23;
  wire and_dcpl_24;
  wire and_dcpl_25;
  wire and_dcpl_26;
  wire and_dcpl_27;
  wire and_dcpl_28;
  wire and_dcpl_29;
  wire and_dcpl_30;
  wire and_dcpl_31;
  wire and_dcpl_32;
  wire and_dcpl_33;
  wire and_dcpl_34;
  wire and_dcpl_35;
  wire and_dcpl_36;
  wire and_dcpl_37;
  wire and_dcpl_38;
  wire and_dcpl_39;
  wire and_dcpl_40;
  wire and_dcpl_41;
  wire and_dcpl_42;
  wire and_dcpl_43;
  wire and_dcpl_44;
  wire and_dcpl_45;
  wire and_dcpl_46;
  wire and_dcpl_47;
  wire and_dcpl_48;
  wire and_dcpl_49;
  wire and_dcpl_50;
  wire and_dcpl_51;
  wire and_dcpl_52;
  wire and_dcpl_53;
  wire and_dcpl_54;
  wire and_dcpl_55;
  wire and_dcpl_56;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire and_dcpl_59;
  wire and_dcpl_60;
  wire and_dcpl_61;
  wire and_dcpl_62;
  wire and_dcpl_63;
  wire and_dcpl_64;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_dcpl_67;
  wire and_dcpl_68;
  wire and_dcpl_69;
  wire and_dcpl_70;
  wire and_dcpl_71;
  wire and_dcpl_72;
  wire and_dcpl_73;
  wire and_dcpl_74;
  wire and_dcpl_75;
  wire and_dcpl_76;
  wire and_dcpl_77;
  wire and_dcpl_78;
  wire and_dcpl_79;
  wire and_dcpl_80;
  wire and_dcpl_81;
  wire and_dcpl_82;
  wire and_dcpl_83;
  wire and_dcpl_84;
  wire and_dcpl_85;
  wire and_dcpl_86;
  wire and_dcpl_87;
  wire and_dcpl_88;
  wire and_dcpl_89;
  wire and_dcpl_90;
  wire and_dcpl_91;
  wire and_dcpl_92;
  wire and_dcpl_93;
  wire and_dcpl_94;
  wire and_dcpl_95;
  wire and_dcpl_96;
  wire and_dcpl_97;
  wire and_dcpl_98;
  wire and_dcpl_99;
  wire and_dcpl_100;
  wire and_dcpl_101;
  wire and_dcpl_102;
  wire and_dcpl_103;
  wire and_dcpl_104;
  wire and_dcpl_105;
  wire and_dcpl_106;
  wire and_dcpl_107;
  wire and_dcpl_108;
  wire and_dcpl_109;
  wire and_dcpl_110;
  wire and_dcpl_111;
  wire and_dcpl_112;
  wire and_dcpl_113;
  wire and_dcpl_114;
  wire and_dcpl_115;
  wire and_dcpl_116;
  wire and_dcpl_117;
  wire and_dcpl_118;
  wire and_dcpl_119;
  wire and_dcpl_120;
  wire and_dcpl_121;
  wire and_dcpl_122;
  wire and_dcpl_123;
  wire and_dcpl_124;
  wire and_dcpl_125;
  wire and_dcpl_126;
  wire and_dcpl_127;
  wire and_dcpl_128;
  wire and_dcpl_129;
  wire and_dcpl_130;
  wire and_dcpl_131;
  wire and_dcpl_132;
  wire and_dcpl_133;
  wire and_dcpl_134;
  wire and_dcpl_135;
  wire and_dcpl_136;
  wire and_dcpl_137;
  wire and_dcpl_138;
  wire and_dcpl_139;
  wire and_dcpl_140;
  wire and_dcpl_141;
  wire and_dcpl_142;
  wire and_dcpl_143;
  wire and_dcpl_144;
  wire and_dcpl_145;
  wire and_dcpl_146;
  wire and_dcpl_147;
  wire and_dcpl_148;
  wire and_dcpl_149;
  wire and_dcpl_150;
  wire and_dcpl_151;
  wire and_dcpl_152;
  wire and_dcpl_153;
  wire and_dcpl_154;
  wire and_dcpl_155;
  wire and_dcpl_156;
  wire and_dcpl_157;
  wire and_dcpl_158;
  wire and_dcpl_159;
  wire and_dcpl_160;
  wire and_dcpl_161;
  wire and_dcpl_162;
  wire and_dcpl_163;
  wire and_dcpl_164;
  wire and_dcpl_165;
  wire and_dcpl_166;
  wire and_dcpl_167;
  wire and_dcpl_168;
  wire and_dcpl_169;
  wire and_dcpl_170;
  wire and_dcpl_171;
  wire and_dcpl_172;
  wire and_dcpl_173;
  wire and_dcpl_174;
  wire and_dcpl_175;
  wire mux_tmp_14;
  wire mux_tmp_15;
  wire and_dcpl_178;
  wire and_dcpl_181;
  wire and_dcpl_187;
  wire and_tmp_1;
  wire mux_tmp_19;
  wire mux_tmp_20;
  wire and_dcpl_188;
  wire and_dcpl_189;
  wire and_dcpl_192;
  wire and_dcpl_195;
  wire or_dcpl_17;
  wire and_dcpl_200;
  reg STORE_OUTPUT_INNER_LOOP_stage_0;
  reg STORE_OUTPUT_INNER_LOOP_stage_0_2;
  reg exit_STORE_OUTPUT_INNER_LOOP_sva_st_1;
  reg [4063:0] reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd;
  reg reg_output_ready_channel_Push_mioi_oswt_cse;
  reg reg_dma_write_chnl_Push_mioi_oswt_cse;
  wire or_15_cse;
  wire or_17_cse;
  wire and_184_rmff;
  wire and_187_rmff;
  reg [31:0] offset_lpi_2;
  reg [24:0] STORE_MAIN_LOOP_s_31_7_sva;
  wire [6:0] STORE_MAIN_LOOP_len_qr_6_0_lpi_2_dfm_1;
  reg [15:0] STORE_OUTPUT_INNER_LOOP_i_sva;
  wire and_dcpl_209;
  wire [31:0] z_out;
  wire [32:0] nl_z_out;
  wire and_dcpl_210;
  wire and_dcpl_211;
  wire and_dcpl_215;
  wire and_dcpl_216;
  wire and_dcpl_217;
  wire and_dcpl_218;
  wire and_dcpl_220;
  wire and_dcpl_221;
  wire and_dcpl_223;
  wire and_dcpl_225;
  wire and_dcpl_227;
  wire and_dcpl_229;
  wire and_dcpl_239;
  wire [24:0] z_out_2;
  wire [25:0] nl_z_out_2;
  reg [63:0] conf_info_crt_2_sva;
  reg [31:0] COMPUTE_BATCH_LOOP_b_sva;
  reg [24:0] STORE_MAIN_LOOP_len_qr_31_7_lpi_2_dfm;
  reg [6:0] STORE_MAIN_LOOP_len_qr_6_0_lpi_2_dfm;
  wire acc_done_mx0c1;
  wire STORE_MAIN_LOOP_len_qr_31_7_lpi_2_dfm_mx0c1;
  wire COMPUTE_BATCH_LOOP_or_1_ssc;
  wire z_out_1_32;

  wire[0:0] mux_12_nl;
  wire[0:0] nor_4_nl;
  wire[0:0] and_203_nl;
  wire[31:0] offset_mul_nl;
  wire[63:0] nl_offset_mul_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] mux_26_nl;
  wire[0:0] mux_25_nl;
  wire[0:0] mux_24_nl;
  wire[0:0] STORE_MAIN_LOOP_len_not_4_nl;
  wire[0:0] or_3_nl;
  wire[0:0] and_23_nl;
  wire[6:0] nor_9_nl;
  wire[6:0] mux1h_nl;
  wire[0:0] mux_21_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] or_18_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] or_16_nl;
  wire[31:0] STORE_MAIN_LOOP_mux_4_nl;
  wire[24:0] STORE_MAIN_LOOP_STORE_MAIN_LOOP_and_1_nl;
  wire[0:0] not_77_nl;
  wire[6:0] STORE_MAIN_LOOP_mux_5_nl;
  wire[33:0] acc_1_nl;
  wire[34:0] nl_acc_1_nl;
  wire[31:0] COMPUTE_BATCH_LOOP_mux1h_3_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_or_2_nl;
  wire[24:0] COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_nor_1_nl;
  wire[24:0] COMPUTE_BATCH_LOOP_mux1h_4_nl;
  wire[6:0] COMPUTE_BATCH_LOOP_mux1h_5_nl;
  wire[24:0] STORE_OUTPUT_INNER_LOOP_mux_2_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output;
  assign nl_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output
      = offset_lpi_2;
  wire[24:0] STORE_MAIN_LOOP_len_qif_mux_nl;
  wire [31:0] nl_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_length_rsc_dat_store_output;
  assign STORE_MAIN_LOOP_len_qif_mux_nl = MUX_v_25_2_2(STORE_MAIN_LOOP_s_31_7_sva,
      25'b0000000000000000000000001, z_out_1_32);
  assign nl_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_length_rsc_dat_store_output
      = {STORE_MAIN_LOOP_len_qif_mux_nl , STORE_MAIN_LOOP_len_qr_6_0_lpi_2_dfm_1};
  wire [63:0] nl_softmax_store_output_store_output_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_m_rsc_dat_store_output;
  assign nl_softmax_store_output_store_output_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_m_rsc_dat_store_output
      = {32'b11011110101011011011111011101111 , STORE_MAIN_LOOP_plm_local_data_rsci_q_d};
  wire [0:0] nl_softmax_store_output_store_output_store_output_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  assign nl_softmax_store_output_store_output_store_output_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0
      = ~ done;
  wire [0:0] nl_softmax_store_output_store_output_store_output_fsm_inst_COMPUTE_BATCH_LOOP_C_0_tr0;
  assign nl_softmax_store_output_store_output_store_output_fsm_inst_COMPUTE_BATCH_LOOP_C_0_tr0
      = ~ z_out_1_32;
  wire [0:0] nl_softmax_store_output_store_output_store_output_fsm_inst_STORE_OUTPUT_INNER_LOOP_C_0_tr0;
  assign nl_softmax_store_output_store_output_store_output_fsm_inst_STORE_OUTPUT_INNER_LOOP_C_0_tr0
      = ~(STORE_OUTPUT_INNER_LOOP_stage_0 | STORE_OUTPUT_INNER_LOOP_stage_0_2);
  wire [0:0] nl_softmax_store_output_store_output_store_output_fsm_inst_STORE_MAIN_LOOP_C_130_tr0;
  assign nl_softmax_store_output_store_output_store_output_fsm_inst_STORE_MAIN_LOOP_C_130_tr0
      = ~ z_out_1_32;
  esp_acc_softmax_softmax_store_output_store_output_output_ready_channel_Push_mioi
      softmax_store_output_store_output_output_ready_channel_Push_mioi_inst (
      .clk(clk),
      .rst(rst),
      .output_ready_channel_val(output_ready_channel_val),
      .output_ready_channel_rdy(output_ready_channel_rdy),
      .output_ready_channel_msg(output_ready_channel_msg),
      .store_output_wen(store_output_wen),
      .output_ready_channel_Push_mioi_oswt(reg_output_ready_channel_Push_mioi_oswt_cse),
      .output_ready_channel_Push_mioi_wen_comp(output_ready_channel_Push_mioi_wen_comp),
      .output_ready_channel_Push_mioi_oswt_pff(and_184_rmff)
    );
  esp_acc_softmax_softmax_store_output_store_output_dma_write_ctrl_Push_mioi softmax_store_output_store_output_dma_write_ctrl_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_ctrl_val(dma_write_ctrl_val),
      .dma_write_ctrl_rdy(dma_write_ctrl_rdy),
      .dma_write_ctrl_msg(dma_write_ctrl_msg),
      .store_output_wen(store_output_wen),
      .dma_write_ctrl_Push_mioi_oswt(reg_output_ready_channel_Push_mioi_oswt_cse),
      .dma_write_ctrl_Push_mioi_wen_comp(dma_write_ctrl_Push_mioi_wen_comp),
      .dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output(nl_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat_store_output[31:0]),
      .dma_write_ctrl_Push_mioi_m_length_rsc_dat_store_output(nl_softmax_store_output_store_output_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_length_rsc_dat_store_output[31:0]),
      .dma_write_ctrl_Push_mioi_oswt_pff(and_184_rmff)
    );
  esp_acc_softmax_softmax_store_output_store_output_dma_write_chnl_Push_mioi softmax_store_output_store_output_dma_write_chnl_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_chnl_val(dma_write_chnl_val),
      .dma_write_chnl_rdy(dma_write_chnl_rdy),
      .dma_write_chnl_msg(dma_write_chnl_msg),
      .store_output_wen(store_output_wen),
      .dma_write_chnl_Push_mioi_oswt(reg_dma_write_chnl_Push_mioi_oswt_cse),
      .dma_write_chnl_Push_mioi_wen_comp(dma_write_chnl_Push_mioi_wen_comp),
      .dma_write_chnl_Push_mioi_m_rsc_dat_store_output(nl_softmax_store_output_store_output_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_m_rsc_dat_store_output[63:0]),
      .dma_write_chnl_Push_mioi_oswt_pff(and_187_rmff)
    );
  esp_acc_softmax_softmax_store_output_store_output_plm_out_cnsi softmax_store_output_store_output_plm_out_cnsi_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_dat(plm_out_cns_dat),
      .plm_out_cns_vld(plm_out_cns_vld),
      .plm_out_cns_rdy(plm_out_cns_rdy),
      .store_output_wen(store_output_wen),
      .plm_out_cnsi_oswt(reg_output_ready_channel_Push_mioi_oswt_cse),
      .plm_out_cnsi_wen_comp(plm_out_cnsi_wen_comp),
      .plm_out_cnsi_idat_mxwt(plm_out_cnsi_idat_mxwt)
    );
  esp_acc_softmax_softmax_store_output_store_output_staller softmax_store_output_store_output_staller_inst
      (
      .store_output_wen(store_output_wen),
      .output_ready_channel_Push_mioi_wen_comp(output_ready_channel_Push_mioi_wen_comp),
      .dma_write_ctrl_Push_mioi_wen_comp(dma_write_ctrl_Push_mioi_wen_comp),
      .dma_write_chnl_Push_mioi_wen_comp(dma_write_chnl_Push_mioi_wen_comp),
      .plm_out_cnsi_wen_comp(plm_out_cnsi_wen_comp)
    );
  esp_acc_softmax_softmax_store_output_store_output_store_output_fsm softmax_store_output_store_output_store_output_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .store_output_wen(store_output_wen),
      .fsm_output(fsm_output),
      .WAIT_FOR_CONFIG_LOOP_C_0_tr0(nl_softmax_store_output_store_output_store_output_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0[0:0]),
      .store_output_rlp_C_0_tr0(z_out_1_32),
      .COMPUTE_BATCH_LOOP_C_0_tr0(nl_softmax_store_output_store_output_store_output_fsm_inst_COMPUTE_BATCH_LOOP_C_0_tr0[0:0]),
      .STORE_OUTPUT_INNER_LOOP_C_0_tr0(nl_softmax_store_output_store_output_store_output_fsm_inst_STORE_OUTPUT_INNER_LOOP_C_0_tr0[0:0]),
      .STORE_MAIN_LOOP_C_130_tr0(nl_softmax_store_output_store_output_store_output_fsm_inst_STORE_MAIN_LOOP_C_130_tr0[0:0]),
      .COMPUTE_BATCH_LOOP_C_1_tr0(z_out_1_32)
    );
  assign STORE_MAIN_LOOP_plm_local_data_rsci_clken_d = store_output_wen;
  assign or_15_cse = (fsm_output[1]) | (fsm_output[3]) | (fsm_output[6]);
  assign and_184_rmff = and_dcpl_18 & and_dcpl_53;
  assign and_187_rmff = and_dcpl_181 & and_dcpl_178 & STORE_OUTPUT_INNER_LOOP_stage_0_2
      & (~ exit_STORE_OUTPUT_INNER_LOOP_sva_st_1);
  assign STORE_MAIN_LOOP_len_not_4_nl = ~ z_out_1_32;
  assign STORE_MAIN_LOOP_len_qr_6_0_lpi_2_dfm_1 = MUX_v_7_2_2(7'b0000000, (conf_info_crt_2_sva[6:0]),
      STORE_MAIN_LOOP_len_not_4_nl);
  assign and_dcpl_3 = ~((fsm_output[6]) | (fsm_output[3]));
  assign and_dcpl_5 = ~((fsm_output[5:4]!=2'b00));
  assign and_dcpl_8 = ~((fsm_output[2]) | (fsm_output[0]));
  assign and_dcpl_9 = (fsm_output[3]) & (~ (fsm_output[1]));
  assign and_dcpl_10 = and_dcpl_9 & and_dcpl_8;
  assign and_dcpl_12 = and_dcpl_5 & (fsm_output[7:6]==2'b10);
  assign or_dcpl_1 = (fsm_output[5:4]!=2'b00);
  assign and_dcpl_14 = (fsm_output[2]) & (~ (fsm_output[0]));
  assign and_dcpl_15 = ~((fsm_output[3]) | (fsm_output[1]));
  assign and_dcpl_16 = and_dcpl_15 & and_dcpl_14;
  assign and_dcpl_17 = ~((fsm_output[7:6]!=2'b00));
  assign and_dcpl_18 = and_dcpl_5 & and_dcpl_17;
  assign and_dcpl_19 = and_dcpl_18 & and_dcpl_16;
  assign and_dcpl_20 = (fsm_output[2]) & (fsm_output[0]);
  assign and_dcpl_21 = and_dcpl_15 & and_dcpl_20;
  assign and_dcpl_23 = (~ (fsm_output[3])) & (fsm_output[1]);
  assign and_dcpl_24 = and_dcpl_23 & and_dcpl_14;
  assign and_dcpl_25 = and_dcpl_18 & and_dcpl_24;
  assign and_dcpl_26 = and_dcpl_23 & and_dcpl_20;
  assign and_dcpl_27 = and_dcpl_18 & and_dcpl_26;
  assign and_dcpl_28 = and_dcpl_18 & and_dcpl_10;
  assign and_dcpl_29 = (~ (fsm_output[2])) & (fsm_output[0]);
  assign and_dcpl_30 = and_dcpl_9 & and_dcpl_29;
  assign and_dcpl_31 = and_dcpl_18 & and_dcpl_30;
  assign and_dcpl_32 = (fsm_output[3]) & (fsm_output[1]);
  assign and_dcpl_33 = and_dcpl_32 & and_dcpl_8;
  assign and_dcpl_34 = and_dcpl_18 & and_dcpl_33;
  assign and_dcpl_35 = and_dcpl_32 & and_dcpl_29;
  assign and_dcpl_36 = and_dcpl_18 & and_dcpl_35;
  assign and_dcpl_37 = and_dcpl_9 & and_dcpl_14;
  assign and_dcpl_38 = and_dcpl_18 & and_dcpl_37;
  assign and_dcpl_39 = and_dcpl_9 & and_dcpl_20;
  assign and_dcpl_40 = and_dcpl_18 & and_dcpl_39;
  assign and_dcpl_41 = and_dcpl_32 & and_dcpl_14;
  assign and_dcpl_42 = and_dcpl_18 & and_dcpl_41;
  assign and_dcpl_43 = and_dcpl_32 & and_dcpl_20;
  assign and_dcpl_44 = and_dcpl_18 & and_dcpl_43;
  assign and_dcpl_45 = and_dcpl_15 & and_dcpl_8;
  assign and_dcpl_46 = (fsm_output[5:4]==2'b01);
  assign and_dcpl_47 = and_dcpl_46 & and_dcpl_17;
  assign and_dcpl_48 = and_dcpl_47 & and_dcpl_45;
  assign and_dcpl_49 = and_dcpl_15 & and_dcpl_29;
  assign and_dcpl_50 = and_dcpl_47 & and_dcpl_49;
  assign and_dcpl_51 = and_dcpl_23 & and_dcpl_8;
  assign and_dcpl_52 = and_dcpl_47 & and_dcpl_51;
  assign and_dcpl_53 = and_dcpl_23 & and_dcpl_29;
  assign and_dcpl_54 = and_dcpl_47 & and_dcpl_53;
  assign and_dcpl_55 = and_dcpl_47 & and_dcpl_16;
  assign and_dcpl_56 = and_dcpl_47 & and_dcpl_21;
  assign and_dcpl_57 = and_dcpl_47 & and_dcpl_24;
  assign and_dcpl_58 = and_dcpl_47 & and_dcpl_26;
  assign and_dcpl_59 = and_dcpl_47 & and_dcpl_10;
  assign and_dcpl_60 = and_dcpl_47 & and_dcpl_30;
  assign and_dcpl_61 = and_dcpl_47 & and_dcpl_33;
  assign and_dcpl_62 = and_dcpl_47 & and_dcpl_35;
  assign and_dcpl_63 = and_dcpl_47 & and_dcpl_37;
  assign and_dcpl_64 = and_dcpl_47 & and_dcpl_39;
  assign and_dcpl_65 = and_dcpl_47 & and_dcpl_41;
  assign and_dcpl_66 = and_dcpl_47 & and_dcpl_43;
  assign and_dcpl_67 = (fsm_output[5:4]==2'b10);
  assign and_dcpl_68 = and_dcpl_67 & and_dcpl_17;
  assign and_dcpl_69 = and_dcpl_68 & and_dcpl_45;
  assign and_dcpl_70 = and_dcpl_68 & and_dcpl_49;
  assign and_dcpl_71 = and_dcpl_68 & and_dcpl_51;
  assign and_dcpl_72 = and_dcpl_68 & and_dcpl_53;
  assign and_dcpl_73 = and_dcpl_68 & and_dcpl_16;
  assign and_dcpl_74 = and_dcpl_68 & and_dcpl_21;
  assign and_dcpl_75 = and_dcpl_68 & and_dcpl_24;
  assign and_dcpl_76 = and_dcpl_68 & and_dcpl_26;
  assign and_dcpl_77 = and_dcpl_68 & and_dcpl_10;
  assign and_dcpl_78 = and_dcpl_68 & and_dcpl_30;
  assign and_dcpl_79 = and_dcpl_68 & and_dcpl_33;
  assign and_dcpl_80 = and_dcpl_68 & and_dcpl_35;
  assign and_dcpl_81 = and_dcpl_68 & and_dcpl_37;
  assign and_dcpl_82 = and_dcpl_68 & and_dcpl_39;
  assign and_dcpl_83 = and_dcpl_68 & and_dcpl_41;
  assign and_dcpl_84 = and_dcpl_68 & and_dcpl_43;
  assign and_dcpl_85 = (fsm_output[5:4]==2'b11);
  assign and_dcpl_86 = and_dcpl_85 & and_dcpl_17;
  assign and_dcpl_87 = and_dcpl_86 & and_dcpl_45;
  assign and_dcpl_88 = and_dcpl_86 & and_dcpl_49;
  assign and_dcpl_89 = and_dcpl_86 & and_dcpl_51;
  assign and_dcpl_90 = and_dcpl_86 & and_dcpl_53;
  assign and_dcpl_91 = and_dcpl_86 & and_dcpl_16;
  assign and_dcpl_92 = and_dcpl_86 & and_dcpl_21;
  assign and_dcpl_93 = and_dcpl_86 & and_dcpl_24;
  assign and_dcpl_94 = and_dcpl_86 & and_dcpl_26;
  assign and_dcpl_95 = and_dcpl_86 & and_dcpl_10;
  assign and_dcpl_96 = and_dcpl_86 & and_dcpl_30;
  assign and_dcpl_97 = and_dcpl_86 & and_dcpl_33;
  assign and_dcpl_98 = and_dcpl_86 & and_dcpl_35;
  assign and_dcpl_99 = and_dcpl_86 & and_dcpl_37;
  assign and_dcpl_100 = and_dcpl_86 & and_dcpl_39;
  assign and_dcpl_101 = and_dcpl_86 & and_dcpl_41;
  assign and_dcpl_102 = and_dcpl_86 & and_dcpl_43;
  assign and_dcpl_103 = (fsm_output[7:6]==2'b01);
  assign and_dcpl_104 = and_dcpl_5 & and_dcpl_103;
  assign and_dcpl_105 = and_dcpl_104 & and_dcpl_45;
  assign and_dcpl_106 = and_dcpl_104 & and_dcpl_49;
  assign and_dcpl_107 = and_dcpl_104 & and_dcpl_51;
  assign and_dcpl_108 = and_dcpl_104 & and_dcpl_53;
  assign and_dcpl_109 = and_dcpl_104 & and_dcpl_16;
  assign and_dcpl_110 = and_dcpl_104 & and_dcpl_21;
  assign and_dcpl_111 = and_dcpl_104 & and_dcpl_24;
  assign and_dcpl_112 = and_dcpl_104 & and_dcpl_26;
  assign and_dcpl_113 = and_dcpl_104 & and_dcpl_10;
  assign and_dcpl_114 = and_dcpl_104 & and_dcpl_30;
  assign and_dcpl_115 = and_dcpl_104 & and_dcpl_33;
  assign and_dcpl_116 = and_dcpl_104 & and_dcpl_35;
  assign and_dcpl_117 = and_dcpl_104 & and_dcpl_37;
  assign and_dcpl_118 = and_dcpl_104 & and_dcpl_39;
  assign and_dcpl_119 = and_dcpl_104 & and_dcpl_41;
  assign and_dcpl_120 = and_dcpl_104 & and_dcpl_43;
  assign and_dcpl_121 = and_dcpl_46 & and_dcpl_103;
  assign and_dcpl_122 = and_dcpl_121 & and_dcpl_45;
  assign and_dcpl_123 = and_dcpl_121 & and_dcpl_49;
  assign and_dcpl_124 = and_dcpl_121 & and_dcpl_51;
  assign and_dcpl_125 = and_dcpl_121 & and_dcpl_53;
  assign and_dcpl_126 = and_dcpl_121 & and_dcpl_16;
  assign and_dcpl_127 = and_dcpl_121 & and_dcpl_21;
  assign and_dcpl_128 = and_dcpl_121 & and_dcpl_24;
  assign and_dcpl_129 = and_dcpl_121 & and_dcpl_26;
  assign and_dcpl_130 = and_dcpl_121 & and_dcpl_10;
  assign and_dcpl_131 = and_dcpl_121 & and_dcpl_30;
  assign and_dcpl_132 = and_dcpl_121 & and_dcpl_33;
  assign and_dcpl_133 = and_dcpl_121 & and_dcpl_35;
  assign and_dcpl_134 = and_dcpl_121 & and_dcpl_37;
  assign and_dcpl_135 = and_dcpl_121 & and_dcpl_39;
  assign and_dcpl_136 = and_dcpl_121 & and_dcpl_41;
  assign and_dcpl_137 = and_dcpl_121 & and_dcpl_43;
  assign and_dcpl_138 = and_dcpl_67 & and_dcpl_103;
  assign and_dcpl_139 = and_dcpl_138 & and_dcpl_45;
  assign and_dcpl_140 = and_dcpl_138 & and_dcpl_49;
  assign and_dcpl_141 = and_dcpl_138 & and_dcpl_51;
  assign and_dcpl_142 = and_dcpl_138 & and_dcpl_53;
  assign and_dcpl_143 = and_dcpl_138 & and_dcpl_16;
  assign and_dcpl_144 = and_dcpl_138 & and_dcpl_21;
  assign and_dcpl_145 = and_dcpl_138 & and_dcpl_24;
  assign and_dcpl_146 = and_dcpl_138 & and_dcpl_26;
  assign and_dcpl_147 = and_dcpl_138 & and_dcpl_10;
  assign and_dcpl_148 = and_dcpl_138 & and_dcpl_30;
  assign and_dcpl_149 = and_dcpl_138 & and_dcpl_33;
  assign and_dcpl_150 = and_dcpl_138 & and_dcpl_35;
  assign and_dcpl_151 = and_dcpl_138 & and_dcpl_37;
  assign and_dcpl_152 = and_dcpl_138 & and_dcpl_39;
  assign and_dcpl_153 = and_dcpl_138 & and_dcpl_41;
  assign and_dcpl_154 = and_dcpl_138 & and_dcpl_43;
  assign and_dcpl_155 = and_dcpl_85 & and_dcpl_103;
  assign and_dcpl_156 = and_dcpl_155 & and_dcpl_45;
  assign and_dcpl_157 = and_dcpl_155 & and_dcpl_49;
  assign and_dcpl_158 = and_dcpl_155 & and_dcpl_51;
  assign and_dcpl_159 = and_dcpl_155 & and_dcpl_53;
  assign and_dcpl_160 = and_dcpl_155 & and_dcpl_16;
  assign and_dcpl_161 = and_dcpl_155 & and_dcpl_21;
  assign and_dcpl_162 = and_dcpl_155 & and_dcpl_24;
  assign and_dcpl_163 = and_dcpl_155 & and_dcpl_26;
  assign and_dcpl_164 = and_dcpl_155 & and_dcpl_10;
  assign and_dcpl_165 = and_dcpl_155 & and_dcpl_30;
  assign and_dcpl_166 = and_dcpl_155 & and_dcpl_33;
  assign and_dcpl_167 = and_dcpl_155 & and_dcpl_35;
  assign and_dcpl_168 = and_dcpl_155 & and_dcpl_37;
  assign and_dcpl_169 = and_dcpl_155 & and_dcpl_39;
  assign and_dcpl_170 = and_dcpl_155 & and_dcpl_41;
  assign and_dcpl_171 = and_dcpl_155 & and_dcpl_43;
  assign and_dcpl_172 = and_dcpl_12 & and_dcpl_45;
  assign and_dcpl_173 = and_dcpl_12 & and_dcpl_49;
  assign and_dcpl_174 = and_dcpl_12 & and_dcpl_51;
  assign and_dcpl_175 = and_dcpl_12 & and_dcpl_53;
  assign mux_tmp_14 = MUX_s_1_2_2(and_dcpl_5, or_dcpl_1, fsm_output[7]);
  assign or_17_cse = (fsm_output[3]) | (fsm_output[6]);
  assign mux_tmp_15 = MUX_s_1_2_2(mux_tmp_14, (fsm_output[7]), or_17_cse);
  assign and_dcpl_178 = (fsm_output[2:0]==3'b101);
  assign and_dcpl_181 = and_dcpl_5 & (fsm_output[7]) & and_dcpl_3;
  assign and_dcpl_187 = and_dcpl_12 & and_dcpl_26;
  assign and_tmp_1 = (fsm_output[7]) & or_dcpl_1;
  assign mux_tmp_19 = MUX_s_1_2_2(and_tmp_1, (fsm_output[7]), or_17_cse);
  assign or_3_nl = (fsm_output[2:1]!=2'b00);
  assign mux_tmp_20 = MUX_s_1_2_2(mux_tmp_15, mux_tmp_19, or_3_nl);
  assign and_dcpl_188 = and_dcpl_18 & and_dcpl_49;
  assign and_dcpl_189 = and_dcpl_12 & and_dcpl_24;
  assign and_dcpl_192 = (fsm_output[2:1]==2'b01);
  assign and_dcpl_195 = and_dcpl_5 & (~ (fsm_output[7])) & and_dcpl_3;
  assign or_dcpl_17 = or_dcpl_1 | (fsm_output[7:6]!=2'b00);
  assign and_dcpl_200 = and_dcpl_12 & and_dcpl_21;
  assign acc_done_mx0c1 = and_dcpl_12 & and_dcpl_10;
  assign STORE_MAIN_LOOP_len_qr_31_7_lpi_2_dfm_mx0c1 = and_dcpl_195 & and_dcpl_192
      & (fsm_output[0]) & (~ z_out_1_32);
  assign and_23_nl = and_dcpl_18 & and_dcpl_21;
  assign STORE_MAIN_LOOP_plm_local_data_rsci_d_d = MUX1HOT_v_32_128_2((plm_out_cnsi_idat_mxwt[4095:4064]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[31:0]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[4063:4032]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[63:32]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[4031:4000]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[95:64]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3999:3968]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[127:96]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3967:3936]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[159:128]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3935:3904]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[191:160]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3903:3872]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[223:192]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3871:3840]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[255:224]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3839:3808]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[287:256]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3807:3776]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[319:288]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3775:3744]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[351:320]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3743:3712]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[383:352]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3711:3680]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[415:384]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3679:3648]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[447:416]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3647:3616]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[479:448]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3615:3584]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[511:480]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3583:3552]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[543:512]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3551:3520]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[575:544]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3519:3488]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[607:576]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3487:3456]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[639:608]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3455:3424]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[671:640]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3423:3392]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[703:672]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3391:3360]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[735:704]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3359:3328]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[767:736]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3327:3296]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[799:768]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3295:3264]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[831:800]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3263:3232]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[863:832]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3231:3200]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[895:864]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3199:3168]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[927:896]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3167:3136]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[959:928]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3135:3104]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[991:960]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3103:3072]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1023:992]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3071:3040]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1055:1024]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3039:3008]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1087:1056]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[3007:2976]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1119:1088]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2975:2944]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1151:1120]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2943:2912]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1183:1152]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2911:2880]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1215:1184]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2879:2848]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1247:1216]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2847:2816]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1279:1248]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2815:2784]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1311:1280]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2783:2752]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1343:1312]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2751:2720]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1375:1344]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2719:2688]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1407:1376]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2687:2656]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1439:1408]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2655:2624]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1471:1440]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2623:2592]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1503:1472]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2591:2560]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1535:1504]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2559:2528]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1567:1536]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2527:2496]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1599:1568]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2495:2464]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1631:1600]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2463:2432]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1663:1632]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2431:2400]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1695:1664]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2399:2368]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1727:1696]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2367:2336]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1759:1728]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2335:2304]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1791:1760]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2303:2272]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1823:1792]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2271:2240]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1855:1824]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2239:2208]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1887:1856]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2207:2176]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1919:1888]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2175:2144]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1951:1920]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2143:2112]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[1983:1952]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2111:2080]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2015:1984]), (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2079:2048]),
      (reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd[2047:2016]), {and_dcpl_19 , and_23_nl
      , and_dcpl_25 , and_dcpl_27 , and_dcpl_28 , and_dcpl_31 , and_dcpl_34 , and_dcpl_36
      , and_dcpl_38 , and_dcpl_40 , and_dcpl_42 , and_dcpl_44 , and_dcpl_48 , and_dcpl_50
      , and_dcpl_52 , and_dcpl_54 , and_dcpl_55 , and_dcpl_56 , and_dcpl_57 , and_dcpl_58
      , and_dcpl_59 , and_dcpl_60 , and_dcpl_61 , and_dcpl_62 , and_dcpl_63 , and_dcpl_64
      , and_dcpl_65 , and_dcpl_66 , and_dcpl_69 , and_dcpl_70 , and_dcpl_71 , and_dcpl_72
      , and_dcpl_73 , and_dcpl_74 , and_dcpl_75 , and_dcpl_76 , and_dcpl_77 , and_dcpl_78
      , and_dcpl_79 , and_dcpl_80 , and_dcpl_81 , and_dcpl_82 , and_dcpl_83 , and_dcpl_84
      , and_dcpl_87 , and_dcpl_88 , and_dcpl_89 , and_dcpl_90 , and_dcpl_91 , and_dcpl_92
      , and_dcpl_93 , and_dcpl_94 , and_dcpl_95 , and_dcpl_96 , and_dcpl_97 , and_dcpl_98
      , and_dcpl_99 , and_dcpl_100 , and_dcpl_101 , and_dcpl_102 , and_dcpl_105 ,
      and_dcpl_106 , and_dcpl_107 , and_dcpl_108 , and_dcpl_109 , and_dcpl_110 ,
      and_dcpl_111 , and_dcpl_112 , and_dcpl_113 , and_dcpl_114 , and_dcpl_115 ,
      and_dcpl_116 , and_dcpl_117 , and_dcpl_118 , and_dcpl_119 , and_dcpl_120 ,
      and_dcpl_122 , and_dcpl_123 , and_dcpl_124 , and_dcpl_125 , and_dcpl_126 ,
      and_dcpl_127 , and_dcpl_128 , and_dcpl_129 , and_dcpl_130 , and_dcpl_131 ,
      and_dcpl_132 , and_dcpl_133 , and_dcpl_134 , and_dcpl_135 , and_dcpl_136 ,
      and_dcpl_137 , and_dcpl_139 , and_dcpl_140 , and_dcpl_141 , and_dcpl_142 ,
      and_dcpl_143 , and_dcpl_144 , and_dcpl_145 , and_dcpl_146 , and_dcpl_147 ,
      and_dcpl_148 , and_dcpl_149 , and_dcpl_150 , and_dcpl_151 , and_dcpl_152 ,
      and_dcpl_153 , and_dcpl_154 , and_dcpl_156 , and_dcpl_157 , and_dcpl_158 ,
      and_dcpl_159 , and_dcpl_160 , and_dcpl_161 , and_dcpl_162 , and_dcpl_163 ,
      and_dcpl_164 , and_dcpl_165 , and_dcpl_166 , and_dcpl_167 , and_dcpl_168 ,
      and_dcpl_169 , and_dcpl_170 , and_dcpl_171 , and_dcpl_172 , and_dcpl_173 ,
      and_dcpl_174 , and_dcpl_175});
  assign STORE_MAIN_LOOP_plm_local_data_rsci_radr_d = STORE_OUTPUT_INNER_LOOP_i_sva[6:0];
  assign mux1h_nl = MUX1HOT_v_7_126_2(7'b0000001, 7'b1111110, 7'b0000010, 7'b1111101,
      7'b0000011, 7'b1111100, 7'b0000100, 7'b1111011, 7'b0000101, 7'b1111010, 7'b0000110,
      7'b1111001, 7'b0000111, 7'b1111000, 7'b0001000, 7'b1110111, 7'b0001001, 7'b1110110,
      7'b0001010, 7'b1110101, 7'b0001011, 7'b1110100, 7'b0001100, 7'b1110011, 7'b0001101,
      7'b1110010, 7'b0001110, 7'b1110001, 7'b0001111, 7'b1110000, 7'b0010000, 7'b1101111,
      7'b0010001, 7'b1101110, 7'b0010010, 7'b1101101, 7'b0010011, 7'b1101100, 7'b0010100,
      7'b1101011, 7'b0010101, 7'b1101010, 7'b0010110, 7'b1101001, 7'b0010111, 7'b1101000,
      7'b0011000, 7'b1100111, 7'b0011001, 7'b1100110, 7'b0011010, 7'b1100101, 7'b0011011,
      7'b1100100, 7'b0011100, 7'b1100011, 7'b0011101, 7'b1100010, 7'b0011110, 7'b1100001,
      7'b0011111, 7'b1100000, 7'b0100000, 7'b1011111, 7'b0100001, 7'b1011110, 7'b0100010,
      7'b1011101, 7'b0100011, 7'b1011100, 7'b0100100, 7'b1011011, 7'b0100101, 7'b1011010,
      7'b0100110, 7'b1011001, 7'b0100111, 7'b1011000, 7'b0101000, 7'b1010111, 7'b0101001,
      7'b1010110, 7'b0101010, 7'b1010101, 7'b0101011, 7'b1010100, 7'b0101100, 7'b1010011,
      7'b0101101, 7'b1010010, 7'b0101110, 7'b1010001, 7'b0101111, 7'b1010000, 7'b0110000,
      7'b1001111, 7'b0110001, 7'b1001110, 7'b0110010, 7'b1001101, 7'b0110011, 7'b1001100,
      7'b0110100, 7'b1001011, 7'b0110101, 7'b1001010, 7'b0110110, 7'b1001001, 7'b0110111,
      7'b1001000, 7'b0111000, 7'b1000111, 7'b0111001, 7'b1000110, 7'b0111010, 7'b1000101,
      7'b0111011, 7'b1000100, 7'b0111100, 7'b1000011, 7'b0111101, 7'b1000010, 7'b0111110,
      7'b1000001, 7'b0111111, 7'b1000000, {and_dcpl_25 , and_dcpl_27 , and_dcpl_28
      , and_dcpl_31 , and_dcpl_34 , and_dcpl_36 , and_dcpl_38 , and_dcpl_40 , and_dcpl_42
      , and_dcpl_44 , and_dcpl_48 , and_dcpl_50 , and_dcpl_52 , and_dcpl_54 , and_dcpl_55
      , and_dcpl_56 , and_dcpl_57 , and_dcpl_58 , and_dcpl_59 , and_dcpl_60 , and_dcpl_61
      , and_dcpl_62 , and_dcpl_63 , and_dcpl_64 , and_dcpl_65 , and_dcpl_66 , and_dcpl_69
      , and_dcpl_70 , and_dcpl_71 , and_dcpl_72 , and_dcpl_73 , and_dcpl_74 , and_dcpl_75
      , and_dcpl_76 , and_dcpl_77 , and_dcpl_78 , and_dcpl_79 , and_dcpl_80 , and_dcpl_81
      , and_dcpl_82 , and_dcpl_83 , and_dcpl_84 , and_dcpl_87 , and_dcpl_88 , and_dcpl_89
      , and_dcpl_90 , and_dcpl_91 , and_dcpl_92 , and_dcpl_93 , and_dcpl_94 , and_dcpl_95
      , and_dcpl_96 , and_dcpl_97 , and_dcpl_98 , and_dcpl_99 , and_dcpl_100 , and_dcpl_101
      , and_dcpl_102 , and_dcpl_105 , and_dcpl_106 , and_dcpl_107 , and_dcpl_108
      , and_dcpl_109 , and_dcpl_110 , and_dcpl_111 , and_dcpl_112 , and_dcpl_113
      , and_dcpl_114 , and_dcpl_115 , and_dcpl_116 , and_dcpl_117 , and_dcpl_118
      , and_dcpl_119 , and_dcpl_120 , and_dcpl_122 , and_dcpl_123 , and_dcpl_124
      , and_dcpl_125 , and_dcpl_126 , and_dcpl_127 , and_dcpl_128 , and_dcpl_129
      , and_dcpl_130 , and_dcpl_131 , and_dcpl_132 , and_dcpl_133 , and_dcpl_134
      , and_dcpl_135 , and_dcpl_136 , and_dcpl_137 , and_dcpl_139 , and_dcpl_140
      , and_dcpl_141 , and_dcpl_142 , and_dcpl_143 , and_dcpl_144 , and_dcpl_145
      , and_dcpl_146 , and_dcpl_147 , and_dcpl_148 , and_dcpl_149 , and_dcpl_150
      , and_dcpl_151 , and_dcpl_152 , and_dcpl_153 , and_dcpl_154 , and_dcpl_156
      , and_dcpl_157 , and_dcpl_158 , and_dcpl_159 , and_dcpl_160 , and_dcpl_161
      , and_dcpl_162 , and_dcpl_163 , and_dcpl_164 , and_dcpl_165 , and_dcpl_166
      , and_dcpl_167 , and_dcpl_168 , and_dcpl_169 , and_dcpl_170 , and_dcpl_171
      , and_dcpl_172 , and_dcpl_173 , and_dcpl_174 , and_dcpl_175});
  assign or_18_nl = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[6]);
  assign mux_20_nl = MUX_s_1_2_2(mux_tmp_14, (fsm_output[7]), or_18_nl);
  assign or_16_nl = (fsm_output[7]) | and_dcpl_5;
  assign mux_16_nl = MUX_s_1_2_2(or_16_nl, (fsm_output[7]), or_15_cse);
  assign mux_19_nl = MUX_s_1_2_2(mux_tmp_15, mux_16_nl, fsm_output[2]);
  assign mux_21_nl = MUX_s_1_2_2(mux_20_nl, mux_19_nl, fsm_output[0]);
  assign nor_9_nl = ~(MUX_v_7_2_2(mux1h_nl, 7'b1111111, mux_21_nl));
  assign STORE_MAIN_LOOP_plm_local_data_rsci_wadr_d = MUX_v_7_2_2(nor_9_nl, 7'b1111111,
      and_dcpl_19);
  assign STORE_MAIN_LOOP_plm_local_data_rsci_we_d_pff = (or_dcpl_1 | (fsm_output[6])
      | (fsm_output[3]) | (fsm_output[2])) ^ (fsm_output[7]);
  assign STORE_MAIN_LOOP_plm_local_data_rsci_readA_r_ram_ir_internal_RMASK_B_d =
      and_dcpl_181 & and_dcpl_178 & STORE_OUTPUT_INNER_LOOP_stage_0 & z_out_1_32;
  assign and_dcpl_209 = and_dcpl_3 & and_dcpl_5 & (fsm_output[7]) & (fsm_output[2])
      & (fsm_output[1]) & (fsm_output[0]);
  assign and_dcpl_210 = (fsm_output[1:0]==2'b01);
  assign and_dcpl_211 = ~((fsm_output[7]) | (fsm_output[2]));
  assign and_dcpl_215 = (fsm_output[6:3]==4'b0000);
  assign and_dcpl_216 = and_dcpl_215 & and_dcpl_211 & and_dcpl_210;
  assign and_dcpl_217 = (fsm_output[1:0]==2'b11);
  assign and_dcpl_218 = (fsm_output[7]) & (fsm_output[2]);
  assign and_dcpl_220 = and_dcpl_215 & and_dcpl_218 & and_dcpl_217;
  assign and_dcpl_221 = (fsm_output[1:0]==2'b10);
  assign and_dcpl_223 = and_dcpl_215 & and_dcpl_211 & and_dcpl_221;
  assign and_dcpl_225 = and_dcpl_215 & and_dcpl_218 & and_dcpl_221;
  assign and_dcpl_227 = and_dcpl_215 & and_dcpl_211 & and_dcpl_217;
  assign and_dcpl_229 = and_dcpl_215 & and_dcpl_218 & and_dcpl_210;
  assign and_dcpl_239 = and_dcpl_3 & and_dcpl_5 & (fsm_output[7]) & (fsm_output[2])
      & (fsm_output[1]) & (~ (fsm_output[0]));
  assign COMPUTE_BATCH_LOOP_or_1_ssc = and_dcpl_216 | and_dcpl_223 | and_dcpl_225;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      acc_done <= 1'b0;
    end
    else if ( store_output_wen & ((mux_12_nl & and_dcpl_5 & and_dcpl_3 & (fsm_output[0])
        & (~ z_out_1_32)) | acc_done_mx0c1) ) begin
      acc_done <= ~ acc_done_mx0c1;
    end
  end
  always @(posedge clk) begin
    if ( store_output_wen ) begin
      conf_info_crt_2_sva <= MUX_v_64_2_2(conf_info_crt_2_sva, conf_info, mux_tmp_20);
      offset_lpi_2 <= MUX1HOT_v_32_3_2(offset_mul_nl, z_out, offset_lpi_2, {and_dcpl_188
          , and_dcpl_189 , (~ mux_27_nl)});
      STORE_OUTPUT_INNER_LOOP_i_sva <= MUX_v_16_2_2(16'b0000000000000000, (z_out_2[15:0]),
          and_dcpl_200);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_output_ready_channel_Push_mioi_oswt_cse <= 1'b0;
      reg_dma_write_chnl_Push_mioi_oswt_cse <= 1'b0;
      exit_STORE_OUTPUT_INNER_LOOP_sva_st_1 <= 1'b0;
      STORE_OUTPUT_INNER_LOOP_stage_0 <= 1'b0;
      STORE_OUTPUT_INNER_LOOP_stage_0_2 <= 1'b0;
    end
    else if ( store_output_wen ) begin
      reg_output_ready_channel_Push_mioi_oswt_cse <= and_184_rmff;
      reg_dma_write_chnl_Push_mioi_oswt_cse <= and_187_rmff;
      exit_STORE_OUTPUT_INNER_LOOP_sva_st_1 <= ~ z_out_1_32;
      STORE_OUTPUT_INNER_LOOP_stage_0 <= ~((~(STORE_OUTPUT_INNER_LOOP_stage_0 & z_out_1_32))
          & and_dcpl_200);
      STORE_OUTPUT_INNER_LOOP_stage_0_2 <= STORE_OUTPUT_INNER_LOOP_stage_0 & and_dcpl_200;
    end
  end
  always @(posedge clk) begin
    if ( store_output_wen & (and_dcpl_188 | and_dcpl_187) ) begin
      COMPUTE_BATCH_LOOP_b_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          z_out, and_dcpl_187);
    end
  end
  always @(posedge clk) begin
    if ( store_output_wen & ((and_dcpl_18 & and_dcpl_51) | and_dcpl_189) ) begin
      STORE_MAIN_LOOP_s_31_7_sva <= MUX_v_25_2_2((conf_info_crt_2_sva[31:7]), z_out_2,
          and_dcpl_189);
    end
  end
  always @(posedge clk) begin
    if ( store_output_wen & ((and_dcpl_195 & and_dcpl_192 & (fsm_output[0]) & z_out_1_32)
        | STORE_MAIN_LOOP_len_qr_31_7_lpi_2_dfm_mx0c1) ) begin
      STORE_MAIN_LOOP_len_qr_31_7_lpi_2_dfm <= MUX_v_25_2_2(25'b0000000000000000000000001,
          STORE_MAIN_LOOP_s_31_7_sva, STORE_MAIN_LOOP_len_qr_31_7_lpi_2_dfm_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( store_output_wen & (~(or_dcpl_17 | (fsm_output[3:0]!=4'b0011))) ) begin
      STORE_MAIN_LOOP_len_qr_6_0_lpi_2_dfm <= STORE_MAIN_LOOP_len_qr_6_0_lpi_2_dfm_1;
    end
  end
  always @(posedge clk) begin
    if ( store_output_wen & (~(or_dcpl_17 | (fsm_output[3:0]!=4'b0100))) ) begin
      reg_STORE_MAIN_LOOP_plm_local_data_asd_ftd <= plm_out_cnsi_idat_mxwt[4063:0];
    end
  end
  assign nor_4_nl = ~((fsm_output[1]) | (fsm_output[7]));
  assign and_203_nl = (fsm_output[1]) & (fsm_output[7]);
  assign mux_12_nl = MUX_s_1_2_2(nor_4_nl, and_203_nl, fsm_output[2]);
  assign nl_offset_mul_nl = (conf_info[31:0]) * (conf_info[63:32]);
  assign offset_mul_nl = nl_offset_mul_nl[31:0];
  assign mux_25_nl = MUX_s_1_2_2(mux_tmp_15, mux_tmp_19, fsm_output[1]);
  assign mux_24_nl = MUX_s_1_2_2(and_tmp_1, (fsm_output[7]), or_15_cse);
  assign mux_26_nl = MUX_s_1_2_2(mux_25_nl, mux_24_nl, fsm_output[2]);
  assign mux_27_nl = MUX_s_1_2_2(mux_26_nl, mux_tmp_20, fsm_output[0]);
  assign STORE_MAIN_LOOP_mux_4_nl = MUX_v_32_2_2(offset_lpi_2, COMPUTE_BATCH_LOOP_b_sva,
      and_dcpl_209);
  assign not_77_nl = ~ and_dcpl_209;
  assign STORE_MAIN_LOOP_STORE_MAIN_LOOP_and_1_nl = MUX_v_25_2_2(25'b0000000000000000000000000,
      STORE_MAIN_LOOP_len_qr_31_7_lpi_2_dfm, not_77_nl);
  assign STORE_MAIN_LOOP_mux_5_nl = MUX_v_7_2_2(STORE_MAIN_LOOP_len_qr_6_0_lpi_2_dfm,
      7'b0000001, and_dcpl_209);
  assign nl_z_out = STORE_MAIN_LOOP_mux_4_nl + ({STORE_MAIN_LOOP_STORE_MAIN_LOOP_and_1_nl
      , STORE_MAIN_LOOP_mux_5_nl});
  assign z_out = nl_z_out[31:0];
  assign COMPUTE_BATCH_LOOP_mux1h_3_nl = MUX1HOT_v_32_6_2((~ (conf_info[63:32])),
      z_out, (~ (conf_info_crt_2_sva[31:0])), ({(~ z_out_2) , (~ (conf_info_crt_2_sva[6:0]))}),
      32'b00000000000000000000000010000001, ({16'b0000000000000000 , STORE_OUTPUT_INNER_LOOP_i_sva}),
      {and_dcpl_216 , and_dcpl_220 , and_dcpl_223 , and_dcpl_225 , and_dcpl_227 ,
      and_dcpl_229});
  assign COMPUTE_BATCH_LOOP_or_2_nl = (~(and_dcpl_216 | and_dcpl_223 | and_dcpl_225
      | and_dcpl_227)) | and_dcpl_220 | and_dcpl_229;
  assign COMPUTE_BATCH_LOOP_mux1h_4_nl = MUX1HOT_v_25_3_2((conf_info_crt_2_sva[63:39]),
      STORE_MAIN_LOOP_s_31_7_sva, STORE_MAIN_LOOP_len_qr_31_7_lpi_2_dfm, {and_dcpl_220
      , and_dcpl_227 , and_dcpl_229});
  assign COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_nor_1_nl = ~(MUX_v_25_2_2(COMPUTE_BATCH_LOOP_mux1h_4_nl,
      25'b1111111111111111111111111, COMPUTE_BATCH_LOOP_or_1_ssc));
  assign COMPUTE_BATCH_LOOP_mux1h_5_nl = MUX1HOT_v_7_4_2(7'b0000001, (~ (conf_info_crt_2_sva[38:32])),
      (~ (conf_info_crt_2_sva[6:0])), (~ STORE_MAIN_LOOP_len_qr_6_0_lpi_2_dfm), {COMPUTE_BATCH_LOOP_or_1_ssc
      , and_dcpl_220 , and_dcpl_227 , and_dcpl_229});
  assign nl_acc_1_nl = ({1'b1 , COMPUTE_BATCH_LOOP_mux1h_3_nl , COMPUTE_BATCH_LOOP_or_2_nl})
      + conv_u2u_33_34({COMPUTE_BATCH_LOOP_COMPUTE_BATCH_LOOP_nor_1_nl , COMPUTE_BATCH_LOOP_mux1h_5_nl
      , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[33:0];
  assign z_out_1_32 = readslicef_34_1_33(acc_1_nl);
  assign STORE_OUTPUT_INNER_LOOP_mux_2_nl = MUX_v_25_2_2(({9'b000000000 , STORE_OUTPUT_INNER_LOOP_i_sva}),
      STORE_MAIN_LOOP_s_31_7_sva, and_dcpl_239);
  assign nl_z_out_2 = STORE_OUTPUT_INNER_LOOP_mux_2_nl + conv_s2u_2_25({and_dcpl_239
      , 1'b1});
  assign z_out_2 = nl_z_out_2[24:0];

  function automatic [24:0] MUX1HOT_v_25_3_2;
    input [24:0] input_2;
    input [24:0] input_1;
    input [24:0] input_0;
    input [2:0] sel;
    reg [24:0] result;
  begin
    result = input_0 & {25{sel[0]}};
    result = result | ( input_1 & {25{sel[1]}});
    result = result | ( input_2 & {25{sel[2]}});
    MUX1HOT_v_25_3_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_128_2;
    input [31:0] input_127;
    input [31:0] input_126;
    input [31:0] input_125;
    input [31:0] input_124;
    input [31:0] input_123;
    input [31:0] input_122;
    input [31:0] input_121;
    input [31:0] input_120;
    input [31:0] input_119;
    input [31:0] input_118;
    input [31:0] input_117;
    input [31:0] input_116;
    input [31:0] input_115;
    input [31:0] input_114;
    input [31:0] input_113;
    input [31:0] input_112;
    input [31:0] input_111;
    input [31:0] input_110;
    input [31:0] input_109;
    input [31:0] input_108;
    input [31:0] input_107;
    input [31:0] input_106;
    input [31:0] input_105;
    input [31:0] input_104;
    input [31:0] input_103;
    input [31:0] input_102;
    input [31:0] input_101;
    input [31:0] input_100;
    input [31:0] input_99;
    input [31:0] input_98;
    input [31:0] input_97;
    input [31:0] input_96;
    input [31:0] input_95;
    input [31:0] input_94;
    input [31:0] input_93;
    input [31:0] input_92;
    input [31:0] input_91;
    input [31:0] input_90;
    input [31:0] input_89;
    input [31:0] input_88;
    input [31:0] input_87;
    input [31:0] input_86;
    input [31:0] input_85;
    input [31:0] input_84;
    input [31:0] input_83;
    input [31:0] input_82;
    input [31:0] input_81;
    input [31:0] input_80;
    input [31:0] input_79;
    input [31:0] input_78;
    input [31:0] input_77;
    input [31:0] input_76;
    input [31:0] input_75;
    input [31:0] input_74;
    input [31:0] input_73;
    input [31:0] input_72;
    input [31:0] input_71;
    input [31:0] input_70;
    input [31:0] input_69;
    input [31:0] input_68;
    input [31:0] input_67;
    input [31:0] input_66;
    input [31:0] input_65;
    input [31:0] input_64;
    input [31:0] input_63;
    input [31:0] input_62;
    input [31:0] input_61;
    input [31:0] input_60;
    input [31:0] input_59;
    input [31:0] input_58;
    input [31:0] input_57;
    input [31:0] input_56;
    input [31:0] input_55;
    input [31:0] input_54;
    input [31:0] input_53;
    input [31:0] input_52;
    input [31:0] input_51;
    input [31:0] input_50;
    input [31:0] input_49;
    input [31:0] input_48;
    input [31:0] input_47;
    input [31:0] input_46;
    input [31:0] input_45;
    input [31:0] input_44;
    input [31:0] input_43;
    input [31:0] input_42;
    input [31:0] input_41;
    input [31:0] input_40;
    input [31:0] input_39;
    input [31:0] input_38;
    input [31:0] input_37;
    input [31:0] input_36;
    input [31:0] input_35;
    input [31:0] input_34;
    input [31:0] input_33;
    input [31:0] input_32;
    input [31:0] input_31;
    input [31:0] input_30;
    input [31:0] input_29;
    input [31:0] input_28;
    input [31:0] input_27;
    input [31:0] input_26;
    input [31:0] input_25;
    input [31:0] input_24;
    input [31:0] input_23;
    input [31:0] input_22;
    input [31:0] input_21;
    input [31:0] input_20;
    input [31:0] input_19;
    input [31:0] input_18;
    input [31:0] input_17;
    input [31:0] input_16;
    input [31:0] input_15;
    input [31:0] input_14;
    input [31:0] input_13;
    input [31:0] input_12;
    input [31:0] input_11;
    input [31:0] input_10;
    input [31:0] input_9;
    input [31:0] input_8;
    input [31:0] input_7;
    input [31:0] input_6;
    input [31:0] input_5;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [127:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    result = result | ( input_5 & {32{sel[5]}});
    result = result | ( input_6 & {32{sel[6]}});
    result = result | ( input_7 & {32{sel[7]}});
    result = result | ( input_8 & {32{sel[8]}});
    result = result | ( input_9 & {32{sel[9]}});
    result = result | ( input_10 & {32{sel[10]}});
    result = result | ( input_11 & {32{sel[11]}});
    result = result | ( input_12 & {32{sel[12]}});
    result = result | ( input_13 & {32{sel[13]}});
    result = result | ( input_14 & {32{sel[14]}});
    result = result | ( input_15 & {32{sel[15]}});
    result = result | ( input_16 & {32{sel[16]}});
    result = result | ( input_17 & {32{sel[17]}});
    result = result | ( input_18 & {32{sel[18]}});
    result = result | ( input_19 & {32{sel[19]}});
    result = result | ( input_20 & {32{sel[20]}});
    result = result | ( input_21 & {32{sel[21]}});
    result = result | ( input_22 & {32{sel[22]}});
    result = result | ( input_23 & {32{sel[23]}});
    result = result | ( input_24 & {32{sel[24]}});
    result = result | ( input_25 & {32{sel[25]}});
    result = result | ( input_26 & {32{sel[26]}});
    result = result | ( input_27 & {32{sel[27]}});
    result = result | ( input_28 & {32{sel[28]}});
    result = result | ( input_29 & {32{sel[29]}});
    result = result | ( input_30 & {32{sel[30]}});
    result = result | ( input_31 & {32{sel[31]}});
    result = result | ( input_32 & {32{sel[32]}});
    result = result | ( input_33 & {32{sel[33]}});
    result = result | ( input_34 & {32{sel[34]}});
    result = result | ( input_35 & {32{sel[35]}});
    result = result | ( input_36 & {32{sel[36]}});
    result = result | ( input_37 & {32{sel[37]}});
    result = result | ( input_38 & {32{sel[38]}});
    result = result | ( input_39 & {32{sel[39]}});
    result = result | ( input_40 & {32{sel[40]}});
    result = result | ( input_41 & {32{sel[41]}});
    result = result | ( input_42 & {32{sel[42]}});
    result = result | ( input_43 & {32{sel[43]}});
    result = result | ( input_44 & {32{sel[44]}});
    result = result | ( input_45 & {32{sel[45]}});
    result = result | ( input_46 & {32{sel[46]}});
    result = result | ( input_47 & {32{sel[47]}});
    result = result | ( input_48 & {32{sel[48]}});
    result = result | ( input_49 & {32{sel[49]}});
    result = result | ( input_50 & {32{sel[50]}});
    result = result | ( input_51 & {32{sel[51]}});
    result = result | ( input_52 & {32{sel[52]}});
    result = result | ( input_53 & {32{sel[53]}});
    result = result | ( input_54 & {32{sel[54]}});
    result = result | ( input_55 & {32{sel[55]}});
    result = result | ( input_56 & {32{sel[56]}});
    result = result | ( input_57 & {32{sel[57]}});
    result = result | ( input_58 & {32{sel[58]}});
    result = result | ( input_59 & {32{sel[59]}});
    result = result | ( input_60 & {32{sel[60]}});
    result = result | ( input_61 & {32{sel[61]}});
    result = result | ( input_62 & {32{sel[62]}});
    result = result | ( input_63 & {32{sel[63]}});
    result = result | ( input_64 & {32{sel[64]}});
    result = result | ( input_65 & {32{sel[65]}});
    result = result | ( input_66 & {32{sel[66]}});
    result = result | ( input_67 & {32{sel[67]}});
    result = result | ( input_68 & {32{sel[68]}});
    result = result | ( input_69 & {32{sel[69]}});
    result = result | ( input_70 & {32{sel[70]}});
    result = result | ( input_71 & {32{sel[71]}});
    result = result | ( input_72 & {32{sel[72]}});
    result = result | ( input_73 & {32{sel[73]}});
    result = result | ( input_74 & {32{sel[74]}});
    result = result | ( input_75 & {32{sel[75]}});
    result = result | ( input_76 & {32{sel[76]}});
    result = result | ( input_77 & {32{sel[77]}});
    result = result | ( input_78 & {32{sel[78]}});
    result = result | ( input_79 & {32{sel[79]}});
    result = result | ( input_80 & {32{sel[80]}});
    result = result | ( input_81 & {32{sel[81]}});
    result = result | ( input_82 & {32{sel[82]}});
    result = result | ( input_83 & {32{sel[83]}});
    result = result | ( input_84 & {32{sel[84]}});
    result = result | ( input_85 & {32{sel[85]}});
    result = result | ( input_86 & {32{sel[86]}});
    result = result | ( input_87 & {32{sel[87]}});
    result = result | ( input_88 & {32{sel[88]}});
    result = result | ( input_89 & {32{sel[89]}});
    result = result | ( input_90 & {32{sel[90]}});
    result = result | ( input_91 & {32{sel[91]}});
    result = result | ( input_92 & {32{sel[92]}});
    result = result | ( input_93 & {32{sel[93]}});
    result = result | ( input_94 & {32{sel[94]}});
    result = result | ( input_95 & {32{sel[95]}});
    result = result | ( input_96 & {32{sel[96]}});
    result = result | ( input_97 & {32{sel[97]}});
    result = result | ( input_98 & {32{sel[98]}});
    result = result | ( input_99 & {32{sel[99]}});
    result = result | ( input_100 & {32{sel[100]}});
    result = result | ( input_101 & {32{sel[101]}});
    result = result | ( input_102 & {32{sel[102]}});
    result = result | ( input_103 & {32{sel[103]}});
    result = result | ( input_104 & {32{sel[104]}});
    result = result | ( input_105 & {32{sel[105]}});
    result = result | ( input_106 & {32{sel[106]}});
    result = result | ( input_107 & {32{sel[107]}});
    result = result | ( input_108 & {32{sel[108]}});
    result = result | ( input_109 & {32{sel[109]}});
    result = result | ( input_110 & {32{sel[110]}});
    result = result | ( input_111 & {32{sel[111]}});
    result = result | ( input_112 & {32{sel[112]}});
    result = result | ( input_113 & {32{sel[113]}});
    result = result | ( input_114 & {32{sel[114]}});
    result = result | ( input_115 & {32{sel[115]}});
    result = result | ( input_116 & {32{sel[116]}});
    result = result | ( input_117 & {32{sel[117]}});
    result = result | ( input_118 & {32{sel[118]}});
    result = result | ( input_119 & {32{sel[119]}});
    result = result | ( input_120 & {32{sel[120]}});
    result = result | ( input_121 & {32{sel[121]}});
    result = result | ( input_122 & {32{sel[122]}});
    result = result | ( input_123 & {32{sel[123]}});
    result = result | ( input_124 & {32{sel[124]}});
    result = result | ( input_125 & {32{sel[125]}});
    result = result | ( input_126 & {32{sel[126]}});
    result = result | ( input_127 & {32{sel[127]}});
    MUX1HOT_v_32_128_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_6_2;
    input [31:0] input_5;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [5:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    result = result | ( input_5 & {32{sel[5]}});
    MUX1HOT_v_32_6_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_126_2;
    input [6:0] input_125;
    input [6:0] input_124;
    input [6:0] input_123;
    input [6:0] input_122;
    input [6:0] input_121;
    input [6:0] input_120;
    input [6:0] input_119;
    input [6:0] input_118;
    input [6:0] input_117;
    input [6:0] input_116;
    input [6:0] input_115;
    input [6:0] input_114;
    input [6:0] input_113;
    input [6:0] input_112;
    input [6:0] input_111;
    input [6:0] input_110;
    input [6:0] input_109;
    input [6:0] input_108;
    input [6:0] input_107;
    input [6:0] input_106;
    input [6:0] input_105;
    input [6:0] input_104;
    input [6:0] input_103;
    input [6:0] input_102;
    input [6:0] input_101;
    input [6:0] input_100;
    input [6:0] input_99;
    input [6:0] input_98;
    input [6:0] input_97;
    input [6:0] input_96;
    input [6:0] input_95;
    input [6:0] input_94;
    input [6:0] input_93;
    input [6:0] input_92;
    input [6:0] input_91;
    input [6:0] input_90;
    input [6:0] input_89;
    input [6:0] input_88;
    input [6:0] input_87;
    input [6:0] input_86;
    input [6:0] input_85;
    input [6:0] input_84;
    input [6:0] input_83;
    input [6:0] input_82;
    input [6:0] input_81;
    input [6:0] input_80;
    input [6:0] input_79;
    input [6:0] input_78;
    input [6:0] input_77;
    input [6:0] input_76;
    input [6:0] input_75;
    input [6:0] input_74;
    input [6:0] input_73;
    input [6:0] input_72;
    input [6:0] input_71;
    input [6:0] input_70;
    input [6:0] input_69;
    input [6:0] input_68;
    input [6:0] input_67;
    input [6:0] input_66;
    input [6:0] input_65;
    input [6:0] input_64;
    input [6:0] input_63;
    input [6:0] input_62;
    input [6:0] input_61;
    input [6:0] input_60;
    input [6:0] input_59;
    input [6:0] input_58;
    input [6:0] input_57;
    input [6:0] input_56;
    input [6:0] input_55;
    input [6:0] input_54;
    input [6:0] input_53;
    input [6:0] input_52;
    input [6:0] input_51;
    input [6:0] input_50;
    input [6:0] input_49;
    input [6:0] input_48;
    input [6:0] input_47;
    input [6:0] input_46;
    input [6:0] input_45;
    input [6:0] input_44;
    input [6:0] input_43;
    input [6:0] input_42;
    input [6:0] input_41;
    input [6:0] input_40;
    input [6:0] input_39;
    input [6:0] input_38;
    input [6:0] input_37;
    input [6:0] input_36;
    input [6:0] input_35;
    input [6:0] input_34;
    input [6:0] input_33;
    input [6:0] input_32;
    input [6:0] input_31;
    input [6:0] input_30;
    input [6:0] input_29;
    input [6:0] input_28;
    input [6:0] input_27;
    input [6:0] input_26;
    input [6:0] input_25;
    input [6:0] input_24;
    input [6:0] input_23;
    input [6:0] input_22;
    input [6:0] input_21;
    input [6:0] input_20;
    input [6:0] input_19;
    input [6:0] input_18;
    input [6:0] input_17;
    input [6:0] input_16;
    input [6:0] input_15;
    input [6:0] input_14;
    input [6:0] input_13;
    input [6:0] input_12;
    input [6:0] input_11;
    input [6:0] input_10;
    input [6:0] input_9;
    input [6:0] input_8;
    input [6:0] input_7;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [125:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    result = result | ( input_3 & {7{sel[3]}});
    result = result | ( input_4 & {7{sel[4]}});
    result = result | ( input_5 & {7{sel[5]}});
    result = result | ( input_6 & {7{sel[6]}});
    result = result | ( input_7 & {7{sel[7]}});
    result = result | ( input_8 & {7{sel[8]}});
    result = result | ( input_9 & {7{sel[9]}});
    result = result | ( input_10 & {7{sel[10]}});
    result = result | ( input_11 & {7{sel[11]}});
    result = result | ( input_12 & {7{sel[12]}});
    result = result | ( input_13 & {7{sel[13]}});
    result = result | ( input_14 & {7{sel[14]}});
    result = result | ( input_15 & {7{sel[15]}});
    result = result | ( input_16 & {7{sel[16]}});
    result = result | ( input_17 & {7{sel[17]}});
    result = result | ( input_18 & {7{sel[18]}});
    result = result | ( input_19 & {7{sel[19]}});
    result = result | ( input_20 & {7{sel[20]}});
    result = result | ( input_21 & {7{sel[21]}});
    result = result | ( input_22 & {7{sel[22]}});
    result = result | ( input_23 & {7{sel[23]}});
    result = result | ( input_24 & {7{sel[24]}});
    result = result | ( input_25 & {7{sel[25]}});
    result = result | ( input_26 & {7{sel[26]}});
    result = result | ( input_27 & {7{sel[27]}});
    result = result | ( input_28 & {7{sel[28]}});
    result = result | ( input_29 & {7{sel[29]}});
    result = result | ( input_30 & {7{sel[30]}});
    result = result | ( input_31 & {7{sel[31]}});
    result = result | ( input_32 & {7{sel[32]}});
    result = result | ( input_33 & {7{sel[33]}});
    result = result | ( input_34 & {7{sel[34]}});
    result = result | ( input_35 & {7{sel[35]}});
    result = result | ( input_36 & {7{sel[36]}});
    result = result | ( input_37 & {7{sel[37]}});
    result = result | ( input_38 & {7{sel[38]}});
    result = result | ( input_39 & {7{sel[39]}});
    result = result | ( input_40 & {7{sel[40]}});
    result = result | ( input_41 & {7{sel[41]}});
    result = result | ( input_42 & {7{sel[42]}});
    result = result | ( input_43 & {7{sel[43]}});
    result = result | ( input_44 & {7{sel[44]}});
    result = result | ( input_45 & {7{sel[45]}});
    result = result | ( input_46 & {7{sel[46]}});
    result = result | ( input_47 & {7{sel[47]}});
    result = result | ( input_48 & {7{sel[48]}});
    result = result | ( input_49 & {7{sel[49]}});
    result = result | ( input_50 & {7{sel[50]}});
    result = result | ( input_51 & {7{sel[51]}});
    result = result | ( input_52 & {7{sel[52]}});
    result = result | ( input_53 & {7{sel[53]}});
    result = result | ( input_54 & {7{sel[54]}});
    result = result | ( input_55 & {7{sel[55]}});
    result = result | ( input_56 & {7{sel[56]}});
    result = result | ( input_57 & {7{sel[57]}});
    result = result | ( input_58 & {7{sel[58]}});
    result = result | ( input_59 & {7{sel[59]}});
    result = result | ( input_60 & {7{sel[60]}});
    result = result | ( input_61 & {7{sel[61]}});
    result = result | ( input_62 & {7{sel[62]}});
    result = result | ( input_63 & {7{sel[63]}});
    result = result | ( input_64 & {7{sel[64]}});
    result = result | ( input_65 & {7{sel[65]}});
    result = result | ( input_66 & {7{sel[66]}});
    result = result | ( input_67 & {7{sel[67]}});
    result = result | ( input_68 & {7{sel[68]}});
    result = result | ( input_69 & {7{sel[69]}});
    result = result | ( input_70 & {7{sel[70]}});
    result = result | ( input_71 & {7{sel[71]}});
    result = result | ( input_72 & {7{sel[72]}});
    result = result | ( input_73 & {7{sel[73]}});
    result = result | ( input_74 & {7{sel[74]}});
    result = result | ( input_75 & {7{sel[75]}});
    result = result | ( input_76 & {7{sel[76]}});
    result = result | ( input_77 & {7{sel[77]}});
    result = result | ( input_78 & {7{sel[78]}});
    result = result | ( input_79 & {7{sel[79]}});
    result = result | ( input_80 & {7{sel[80]}});
    result = result | ( input_81 & {7{sel[81]}});
    result = result | ( input_82 & {7{sel[82]}});
    result = result | ( input_83 & {7{sel[83]}});
    result = result | ( input_84 & {7{sel[84]}});
    result = result | ( input_85 & {7{sel[85]}});
    result = result | ( input_86 & {7{sel[86]}});
    result = result | ( input_87 & {7{sel[87]}});
    result = result | ( input_88 & {7{sel[88]}});
    result = result | ( input_89 & {7{sel[89]}});
    result = result | ( input_90 & {7{sel[90]}});
    result = result | ( input_91 & {7{sel[91]}});
    result = result | ( input_92 & {7{sel[92]}});
    result = result | ( input_93 & {7{sel[93]}});
    result = result | ( input_94 & {7{sel[94]}});
    result = result | ( input_95 & {7{sel[95]}});
    result = result | ( input_96 & {7{sel[96]}});
    result = result | ( input_97 & {7{sel[97]}});
    result = result | ( input_98 & {7{sel[98]}});
    result = result | ( input_99 & {7{sel[99]}});
    result = result | ( input_100 & {7{sel[100]}});
    result = result | ( input_101 & {7{sel[101]}});
    result = result | ( input_102 & {7{sel[102]}});
    result = result | ( input_103 & {7{sel[103]}});
    result = result | ( input_104 & {7{sel[104]}});
    result = result | ( input_105 & {7{sel[105]}});
    result = result | ( input_106 & {7{sel[106]}});
    result = result | ( input_107 & {7{sel[107]}});
    result = result | ( input_108 & {7{sel[108]}});
    result = result | ( input_109 & {7{sel[109]}});
    result = result | ( input_110 & {7{sel[110]}});
    result = result | ( input_111 & {7{sel[111]}});
    result = result | ( input_112 & {7{sel[112]}});
    result = result | ( input_113 & {7{sel[113]}});
    result = result | ( input_114 & {7{sel[114]}});
    result = result | ( input_115 & {7{sel[115]}});
    result = result | ( input_116 & {7{sel[116]}});
    result = result | ( input_117 & {7{sel[117]}});
    result = result | ( input_118 & {7{sel[118]}});
    result = result | ( input_119 & {7{sel[119]}});
    result = result | ( input_120 & {7{sel[120]}});
    result = result | ( input_121 & {7{sel[121]}});
    result = result | ( input_122 & {7{sel[122]}});
    result = result | ( input_123 & {7{sel[123]}});
    result = result | ( input_124 & {7{sel[124]}});
    result = result | ( input_125 & {7{sel[125]}});
    MUX1HOT_v_7_126_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_4_2;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [3:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    result = result | ( input_3 & {7{sel[3]}});
    MUX1HOT_v_7_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [24:0] MUX_v_25_2_2;
    input [24:0] input_0;
    input [24:0] input_1;
    input [0:0] sel;
    reg [24:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_25_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_34_1_33;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 33;
    readslicef_34_1_33 = tmp[0:0];
  end
  endfunction


  function automatic [24:0] conv_s2u_2_25 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_25 = {{23{vector[1]}}, vector};
  end
  endfunction


  function automatic [33:0] conv_u2u_33_34 ;
    input [32:0]  vector ;
  begin
    conv_u2u_33_34 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel_compute_kernel
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel_compute_kernel (
  clk, rst, conf_info, done, input_ready_channel_val, input_ready_channel_rdy, input_ready_channel_msg,
      output_ready_channel_val, output_ready_channel_rdy, output_ready_channel_msg,
      plm_in_cns_dat, plm_in_cns_vld, plm_in_cns_rdy, plm_out_cns_dat, plm_out_cns_vld,
      plm_out_cns_rdy, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_adra_d, COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_da_d,
      COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d, COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_wea_d,
      COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_adra_d, COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_da_d,
      COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d, COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_wea_d,
      COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_adra_d, COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_da_d,
      COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d, COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_wea_d,
      COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_adra_d, COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_da_d,
      COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d, COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_wea_d,
      COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      CALC_SOFTMAX_LOOP_mul_cmp_b, CALC_SOFTMAX_LOOP_mul_cmp_z, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff
);
  input clk;
  input rst;
  input [63:0] conf_info;
  input done;
  output input_ready_channel_val;
  input input_ready_channel_rdy;
  output input_ready_channel_msg;
  input output_ready_channel_val;
  output output_ready_channel_rdy;
  input output_ready_channel_msg;
  input [4095:0] plm_in_cns_dat;
  input plm_in_cns_vld;
  output plm_in_cns_rdy;
  output [4095:0] plm_out_cns_dat;
  output plm_out_cns_vld;
  input plm_out_cns_rdy;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d;
  output [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d;
  output [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d;
  output [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_adra_d;
  output [2047:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_da_d;
  input [2047:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_wea_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_adra_d;
  output [2047:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_da_d;
  input [2047:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_wea_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_adra_d;
  output [1023:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_da_d;
  input [2047:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_wea_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_adra_d;
  output [1023:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_da_d;
  input [2047:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_wea_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  output [93:0] CALC_SOFTMAX_LOOP_mul_cmp_b;
  input [94:0] CALC_SOFTMAX_LOOP_mul_cmp_z;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff;


  // Interconnect Declarations
  wire compute_kernel_wen;
  wire input_ready_channel_Push_mioi_wen_comp;
  wire output_ready_channel_Pop_mioi_wen_comp;
  wire plm_in_cnsi_wen_comp;
  wire [4095:0] plm_in_cnsi_idat_mxwt;
  wire plm_out_cnsi_wen_comp;
  reg [1023:0] plm_out_cnsi_idat_4095_3072;
  reg [1023:0] plm_out_cnsi_idat_3071_2048;
  reg [1023:0] plm_out_cnsi_idat_2047_1024;
  reg [1023:0] plm_out_cnsi_idat_1023_0;
  wire [5:0] fsm_output;
  wire [7:0] CALC_SOFTMAX_LOOP_acc_1_tmp;
  wire [8:0] nl_CALC_SOFTMAX_LOOP_acc_1_tmp;
  wire [73:0] SUM_EXP_LOOP_acc_1_tmp;
  wire [74:0] nl_SUM_EXP_LOOP_acc_1_tmp;
  wire [7:0] SUM_EXP_LOOP_acc_2_tmp;
  wire [8:0] nl_SUM_EXP_LOOP_acc_2_tmp;
  wire [7:0] CALC_EXP_LOOP_acc_1_tmp;
  wire [8:0] nl_CALC_EXP_LOOP_acc_1_tmp;
  wire or_dcpl_6;
  wire and_dcpl_7;
  wire and_dcpl_13;
  wire and_dcpl_87;
  wire or_dcpl_36;
  wire or_dcpl_41;
  wire not_tmp_75;
  wire and_dcpl_108;
  wire and_dcpl_113;
  wire mux_tmp_35;
  wire and_dcpl_114;
  wire and_dcpl_115;
  wire and_dcpl_118;
  wire or_tmp_47;
  wire and_191_cse;
  wire and_192_cse;
  wire and_239_cse;
  reg exitL_exit_CALC_SOFTMAX_LOOP_sva;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_4_1_1;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_4_0_1;
  wire CALC_SOFTMAX_LOOP_or_tmp_1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_66;
  wire CALC_SOFTMAX_LOOP_equal_tmp_67;
  wire exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_1;
  wire CALC_SOFTMAX_LOOP_and_4_ssc_1;
  wire CALC_SOFTMAX_LOOP_and_5_ssc_1;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_0_mx0;
  wire CALC_EXP_LOOP_and_svs_mx1w2;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_1_mx0;
  reg CALC_SOFTMAX_LOOP_nor_26_itm;
  reg CALC_SOFTMAX_LOOP_nor_28_itm;
  reg CALC_SOFTMAX_LOOP_nor_1_itm;
  reg CALC_SOFTMAX_LOOP_nor_25_itm;
  reg CALC_SOFTMAX_LOOP_nor_14_itm;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_0;
  reg COMPUTE_OUTER_LOOP_asn_6_itm_2;
  reg COMPUTE_OUTER_LOOP_stage_0_3;
  reg CALC_SOFTMAX_LOOP_and_10_itm_2;
  reg COMPUTE_OUTER_LOOP_stage_0;
  reg COMPUTE_OUTER_LOOP_stage_0_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_1;
  reg COMPUTE_OUTER_LOOP_stage_0_2;
  reg COMPUTE_OUTER_LOOP_asn_6_itm_1;
  reg COMPUTE_OUTER_LOOP_stage_0_6;
  reg exit_COMPUTE_OUTER_LOOP_sva_1;
  reg CALC_SOFTMAX_LOOP_asn_itm;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_0;
  reg CALC_SOFTMAX_LOOP_and_10_itm;
  reg CALC_SOFTMAX_LOOP_asn_itm_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_10_1;
  reg CALC_SOFTMAX_LOOP_and_10_itm_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_4_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_4_1;
  reg exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_4;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_1;
  reg exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_3;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_2_1;
  reg exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_2;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_2_0;
  reg CALC_SOFTMAX_LOOP_equal_tmp_10_2;
  reg CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_1;
  reg CALC_SOFTMAX_LOOP_asn_3_itm;
  reg COMPUTE_OUTER_LOOP_stage_0_4;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_0;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_4;
  reg CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_itm_1;
  reg CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm;
  reg CALC_SOFTMAX_LOOP_equal_tmp_15;
  reg CALC_SOFTMAX_LOOP_equal_tmp_14;
  reg CALC_SOFTMAX_LOOP_equal_tmp_20;
  reg CALC_SOFTMAX_LOOP_equal_tmp_16;
  reg CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_3_itm;
  reg CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_3;
  reg COMPUTE_OUTER_LOOP_stage_0_5;
  reg CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_itm;
  reg [6:0] CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0;
  reg [6:0] CALC_SOFTMAX_LOOP_i_7_0_lpi_2_dfm_2_6_0;
  reg CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2;
  wire [4:0] CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0;
  wire CALC_SOFTMAX_LOOP_and_7_tmp;
  wire and_138_m1c;
  wire and_121_m1c;
  wire or_162_tmp;
  reg reg_input_ready_channel_Push_mioi_oswt_cse;
  reg reg_output_ready_channel_Pop_mioi_oswt_cse;
  wire COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_nor_cse;
  wire COMPUTE_OUTER_LOOP_and_cse;
  wire or_8_cse;
  wire COMPUTE_OUTER_LOOP_and_4_cse;
  wire and_163_rmff;
  wire COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_mux_7_rmff;
  wire and_189_rmff;
  wire and_210_rmff;
  wire and_150_rmff;
  wire and_152_rmff;
  wire COMPUTE_OUTER_LOOP_nor_2_seb;
  wire COMPUTE_OUTER_LOOP_nor_1_seb;
  reg CALC_SOFTMAX_LOOP_equal_tmp_32_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_31_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_30_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_29_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_28_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_27_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_26_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_25_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_24_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_23_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_22_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_21_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_20_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_19_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_18_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_17_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_16_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_15_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_14_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_13_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_12_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_11_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_10_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_41_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_40_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_39_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_38_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_37_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_36_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_3_3;
  reg CALC_SOFTMAX_LOOP_equal_tmp_2_3;
  wire CALC_SOFTMAX_LOOP_or_152;
  reg [93:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_2;
  wire [66:0] operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1;
  reg [6:0] CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_6_0;
  reg [6:0] CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0;
  reg [73:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_2_dfm_1;
  reg [73:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_2;
  wire or_414_tmp;
  wire [72:0] operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm;
  wire [93:0] operator_94_21_false_AC_TRN_AC_WRAP_rshift_itm;
  wire [31:0] z_out_1;
  wire [32:0] nl_z_out_1;
  reg [63:0] conf_info_crt_1_sva;
  reg [31:0] COMPUTE_BATCH_LOOP_b_sva;
  reg [24:0] COMPUTE_OUTER_LOOP_s_31_7_sva;
  reg [12:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_normalized_fixed_72_60_sva;
  reg CALC_SOFTMAX_LOOP_equal_tmp_5;
  reg CALC_SOFTMAX_LOOP_equal_tmp_22;
  reg CALC_SOFTMAX_LOOP_equal_tmp_23;
  reg CALC_SOFTMAX_LOOP_equal_tmp_24;
  reg CALC_SOFTMAX_LOOP_equal_tmp_26;
  reg CALC_SOFTMAX_LOOP_equal_tmp_27;
  reg CALC_SOFTMAX_LOOP_equal_tmp_28;
  reg CALC_SOFTMAX_LOOP_equal_tmp_29;
  reg CALC_SOFTMAX_LOOP_equal_tmp_30;
  reg CALC_SOFTMAX_LOOP_equal_tmp_31;
  reg CALC_SOFTMAX_LOOP_equal_tmp_32;
  reg CALC_SOFTMAX_LOOP_equal_tmp_64;
  reg [7:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm;
  wire [8:0] nl_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm;
  reg CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_5_itm;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm;
  reg CALC_SOFTMAX_LOOP_equal_tmp_2_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_2_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_3_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_3_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_4_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_4_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_5_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_6_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_6_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_11_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_11_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_12_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_12_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_13_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_13_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_14_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_14_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_15_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_15_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_16_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_16_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_17_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_17_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_18_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_18_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_19_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_19_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_20_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_20_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_21_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_21_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_22_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_22_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_23_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_23_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_24_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_24_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_25_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_25_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_26_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_26_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_27_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_27_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_28_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_28_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_29_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_29_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_30_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_30_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_31_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_31_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_32_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_32_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_62_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_62_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_63_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_63_2;
  reg CALC_SOFTMAX_LOOP_equal_tmp_64_1;
  reg CALC_SOFTMAX_LOOP_equal_tmp_64_2;
  reg [1023:0] tmp_3_sva_1;
  reg [1023:0] tmp_4_sva_1;
  reg [4:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_itm_1;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_1_itm_1;
  reg [9:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_32_14_11_0_1_itm_1;
  reg [2:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_2_itm_1;
  reg [6:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_3_itm_1;
  reg [6:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_32_14_18_12_itm_1;
  reg CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_3_itm_1;
  reg CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_3_itm_2;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_1;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_2;
  reg CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_3;
  reg [6:0] SUM_EXP_LOOP_i_7_0_lpi_2_6_0;
  wire [6:0] CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_44_mx1w0;
  wire CALC_SOFTMAX_LOOP_equal_tmp_40_mx1w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_39_mx1w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_57_mx1w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_53_mx1w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_51_mx1w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_50_mx1w2;
  wire CALC_SOFTMAX_LOOP_equal_tmp_49_mx1w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_45_mx1w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_43_mx1w2;
  wire CALC_SOFTMAX_LOOP_equal_tmp_42_mx1w2;
  wire CALC_SOFTMAX_LOOP_equal_tmp_38_mx1w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_37_mx1w0;
  wire CALC_SOFTMAX_LOOP_equal_tmp_36_mx1w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_2_mx1w0;
  wire CALC_SOFTMAX_LOOP_equal_tmp_46_mx1w0;
  wire CALC_SOFTMAX_LOOP_equal_tmp_47_mx1w0;
  wire CALC_SOFTMAX_LOOP_equal_tmp_48_mx1w0;
  wire CALC_SOFTMAX_LOOP_equal_tmp_52_mx1w0;
  wire [6:0] CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_6_0_mx1;
  wire CALC_SOFTMAX_LOOP_nor_26_itm_mx1w0;
  wire CALC_SOFTMAX_LOOP_nor_32_itm_mx1w1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_and_4_mx0w0;
  wire COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_and_3_mx0w0;
  wire CALC_SOFTMAX_LOOP_equal_tmp_64_mx0w0;
  wire CALC_SOFTMAX_LOOP_equal_tmp_63_mx0w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_62_mx0w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_61_mx0w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_60_mx0w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_59_mx0w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_58_mx0w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_56_mx0w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_55_mx0w1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_54_mx0w1;
  wire [18:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire signed [19:0] nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire [6:0] libraries_leading_sign_74_0_5d32be77710879fd6707bb2fa0416553bf16_1;
  wire or_173_tmp;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_and_6_rgt;
  wire CALC_SOFTMAX_LOOP_i_and_rgt;
  wire CALC_SOFTMAX_LOOP_i_and_1_rgt;
  wire and_140_rgt;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_and_4_rgt;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_and_3_rgt;
  wire and_615_rgt;
  wire COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_or_5_cse;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_and_cse;
  wire CALC_SOFTMAX_LOOP_and_cse;
  wire CALC_SOFTMAX_LOOP_i_and_4_cse;
  wire CALC_SOFTMAX_LOOP_and_79_cse;
  wire CALC_SOFTMAX_LOOP_and_57_cse;
  wire CALC_SOFTMAX_LOOP_and_88_cse;
  wire COMPUTE_OUTER_LOOP_acc_itm_32_1;
  wire [18:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28;
  wire z_out_32;

  wire[0:0] mux_34_nl;
  wire[0:0] or_78_nl;
  wire[0:0] mux_35_nl;
  wire[0:0] or_82_nl;
  wire[93:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_or_nl;
  wire[0:0] and_247_nl;
  wire[0:0] COMPUTE_OUTER_LOOP_mux_33_nl;
  wire[0:0] COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_mux_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_nl;
  wire[0:0] COMPUTE_OUTER_LOOP_and_16_nl;
  wire[0:0] CALC_EXP_LOOP_i_CALC_EXP_LOOP_i_nor_nl;
  wire[0:0] CALC_EXP_LOOP_i_and_1_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux1h_22_nl;
  wire[0:0] COMPUTE_OUTER_LOOP_s_and_nl;
  wire[0:0] COMPUTE_OUTER_LOOP_s_and_2_nl;
  wire[0:0] COMPUTE_OUTER_LOOP_s_or_nl;
  wire[0:0] or_269_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_14_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_16_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_18_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_20_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_22_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_24_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_26_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_28_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_30_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_32_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_34_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_36_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_38_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_40_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_42_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_44_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_46_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_48_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_50_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_52_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_54_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_56_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_58_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_60_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_62_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_64_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_66_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_68_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_70_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_72_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_74_nl;
  wire[0:0] COMPUTE_OUTER_LOOP_mux_32_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_10_nl;
  wire[0:0] nor_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_41_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_35_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_68_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_4_nl;
  wire[31:0] COMPUTE_BATCH_LOOP_b_mux_nl;
  wire[0:0] softmax_softmax_not_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_and_10_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_164_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_166_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_168_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_170_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux1h_228_nl;
  wire[32:0] COMPUTE_OUTER_LOOP_acc_nl;
  wire[33:0] nl_COMPUTE_OUTER_LOOP_acc_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_183_nl;
  wire[6:0] CALC_SOFTMAX_LOOP_mux_184_nl;
  wire[7:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_nl;
  wire[46:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl;
  wire signed [47:0] nl_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_5_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_6_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_7_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_8_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_9_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_10_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_11_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_12_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_13_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_14_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_15_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_16_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_17_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_18_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_19_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_20_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_21_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_22_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_23_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_24_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_25_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_26_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_27_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_28_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_29_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_30_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_31_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_32_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_33_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_34_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_35_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_36_nl;
  wire[31:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_37_nl;
  wire[0:0] nor_13_nl;
  wire[0:0] or_168_nl;
  wire[0:0] COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_or_1_nl;
  wire[0:0] and_166_nl;
  wire[0:0] COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_and_nl;
  wire[0:0] and_178_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_1_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_2_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_3_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_4_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_5_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_6_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_7_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_8_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_9_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_10_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_11_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_12_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_13_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_14_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_15_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_16_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_17_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_18_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_19_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_20_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_21_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_22_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_23_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_24_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_25_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_26_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_27_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_28_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_29_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_30_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_31_nl;
  wire[0:0] COMPUTE_OUTER_LOOP_and_9_nl;
  wire[0:0] COMPUTE_OUTER_LOOP_and_13_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_32_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_33_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_34_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_35_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_36_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_37_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_38_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_39_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_40_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_41_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_42_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_43_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_44_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_45_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_46_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_47_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_48_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_49_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_50_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_51_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_52_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_53_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_54_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_55_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_56_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_57_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_58_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_59_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_60_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_61_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_62_nl;
  wire[31:0] CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_63_nl;
  wire[0:0] COMPUTE_OUTER_LOOP_and_10_nl;
  wire[0:0] COMPUTE_OUTER_LOOP_and_14_nl;
  wire[33:0] acc_nl;
  wire[34:0] nl_acc_nl;
  wire[31:0] COMPUTE_BATCH_LOOP_mux_4_nl;
  wire[0:0] COMPUTE_BATCH_LOOP_or_1_nl;
  wire[31:0] COMPUTE_BATCH_LOOP_mux_5_nl;
  wire[31:0] COMPUTE_OUTER_LOOP_mux_34_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [72:0] nl_operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg_a = SUM_EXP_LOOP_acc_1_tmp[72:0];
  wire[10:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[9:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl;
  wire [73:0] nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_a;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl
      = MUX_v_10_8_2(10'b1111111101, 10'b1100011001, 10'b1001100100, 10'b0111010000,
      10'b0101010100, 10'b0011101011, 10'b0010010001, 10'b0001000100, ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_normalized_fixed_72_60_sva[12:10]);
  assign nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_s2u_9_11(ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:10])
      + ({1'b1 , ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl});
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_a = {ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , (ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[9:0])
      , 53'b00000000000000000000000000000000000000000000000000000};
  wire[10:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire [20:0] nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:10])
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_2_itm_1
      , 1'b1 , ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_3_itm_1});
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a = {ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , (ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[9:0])};
  wire [4095:0] nl_softmax_compute_kernel_compute_kernel_plm_out_cnsi_inst_plm_out_cnsi_idat;
  assign nl_softmax_compute_kernel_compute_kernel_plm_out_cnsi_inst_plm_out_cnsi_idat
      = {plm_out_cnsi_idat_4095_3072 , plm_out_cnsi_idat_3071_2048 , plm_out_cnsi_idat_2047_1024
      , plm_out_cnsi_idat_1023_0};
  wire [0:0] nl_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  assign nl_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0
      = ~ done;
  wire [0:0] nl_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_inst_COMPUTE_OUTER_LOOP_C_1_tr0;
  assign nl_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_inst_COMPUTE_OUTER_LOOP_C_1_tr0
      = COMPUTE_OUTER_LOOP_stage_0 | COMPUTE_OUTER_LOOP_stage_0_5 | COMPUTE_OUTER_LOOP_stage_0_4
      | COMPUTE_OUTER_LOOP_stage_0_2 | COMPUTE_OUTER_LOOP_stage_0_1 | COMPUTE_OUTER_LOOP_stage_0_3;
  esp_acc_softmax_mgc_shift_l_v5 #(.width_a(32'sd73),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd73)) operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg_a[72:0]),
      .s(libraries_leading_sign_74_0_5d32be77710879fd6707bb2fa0416553bf16_1),
      .z(operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  esp_acc_softmax_mgc_shift_br_v5 #(.width_a(32'sd74),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd94)) operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_a[73:0]),
      .s(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm),
      .z(operator_94_21_false_AC_TRN_AC_WRAP_rshift_itm)
    );
  esp_acc_softmax_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd67)) operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_32_14_18_12_itm_1),
      .z(operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1)
    );
  esp_acc_softmax_leading_sign_74_0  leading_sign_74_0_rg (
      .mantissa(SUM_EXP_LOOP_acc_1_tmp),
      .rtn(libraries_leading_sign_74_0_5d32be77710879fd6707bb2fa0416553bf16_1)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_input_ready_channel_Push_mioi
      softmax_compute_kernel_compute_kernel_input_ready_channel_Push_mioi_inst (
      .clk(clk),
      .rst(rst),
      .input_ready_channel_val(input_ready_channel_val),
      .input_ready_channel_rdy(input_ready_channel_rdy),
      .input_ready_channel_msg(input_ready_channel_msg),
      .compute_kernel_wen(compute_kernel_wen),
      .input_ready_channel_Push_mioi_oswt(reg_input_ready_channel_Push_mioi_oswt_cse),
      .input_ready_channel_Push_mioi_wen_comp(input_ready_channel_Push_mioi_wen_comp),
      .input_ready_channel_Push_mioi_oswt_pff(and_150_rmff)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_output_ready_channel_Pop_mioi
      softmax_compute_kernel_compute_kernel_output_ready_channel_Pop_mioi_inst (
      .clk(clk),
      .rst(rst),
      .output_ready_channel_val(output_ready_channel_val),
      .output_ready_channel_rdy(output_ready_channel_rdy),
      .output_ready_channel_msg(output_ready_channel_msg),
      .compute_kernel_wen(compute_kernel_wen),
      .output_ready_channel_Pop_mioi_oswt(reg_output_ready_channel_Pop_mioi_oswt_cse),
      .output_ready_channel_Pop_mioi_wen_comp(output_ready_channel_Pop_mioi_wen_comp),
      .output_ready_channel_Pop_mioi_oswt_pff(and_152_rmff)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_in_cnsi softmax_compute_kernel_compute_kernel_plm_in_cnsi_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_dat(plm_in_cns_dat),
      .plm_in_cns_vld(plm_in_cns_vld),
      .plm_in_cns_rdy(plm_in_cns_rdy),
      .compute_kernel_wen(compute_kernel_wen),
      .plm_in_cnsi_oswt(reg_input_ready_channel_Push_mioi_oswt_cse),
      .plm_in_cnsi_wen_comp(plm_in_cnsi_wen_comp),
      .plm_in_cnsi_idat_mxwt(plm_in_cnsi_idat_mxwt)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_plm_out_cnsi softmax_compute_kernel_compute_kernel_plm_out_cnsi_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_out_cns_dat(plm_out_cns_dat),
      .plm_out_cns_vld(plm_out_cns_vld),
      .plm_out_cns_rdy(plm_out_cns_rdy),
      .compute_kernel_wen(compute_kernel_wen),
      .plm_out_cnsi_oswt(reg_output_ready_channel_Pop_mioi_oswt_cse),
      .plm_out_cnsi_wen_comp(plm_out_cnsi_wen_comp),
      .plm_out_cnsi_idat(nl_softmax_compute_kernel_compute_kernel_plm_out_cnsi_inst_plm_out_cnsi_idat[4095:0])
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_staller softmax_compute_kernel_compute_kernel_staller_inst
      (
      .compute_kernel_wen(compute_kernel_wen),
      .input_ready_channel_Push_mioi_wen_comp(input_ready_channel_Push_mioi_wen_comp),
      .output_ready_channel_Pop_mioi_wen_comp(output_ready_channel_Pop_mioi_wen_comp),
      .plm_in_cnsi_wen_comp(plm_in_cnsi_wen_comp),
      .plm_out_cnsi_wen_comp(plm_out_cnsi_wen_comp)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel_compute_kernel_fsm softmax_compute_kernel_compute_kernel_compute_kernel_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .compute_kernel_wen(compute_kernel_wen),
      .fsm_output(fsm_output),
      .WAIT_FOR_CONFIG_LOOP_C_0_tr0(nl_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0[0:0]),
      .compute_kernel_rlp_C_0_tr0(z_out_32),
      .COMPUTE_OUTER_LOOP_C_1_tr0(nl_softmax_compute_kernel_compute_kernel_compute_kernel_fsm_inst_COMPUTE_OUTER_LOOP_C_1_tr0[0:0]),
      .COMPUTE_BATCH_LOOP_C_0_tr0(z_out_32)
    );
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d
      = compute_kernel_wen;
  assign and_150_rmff = exitL_exit_CALC_SOFTMAX_LOOP_sva & COMPUTE_OUTER_LOOP_acc_itm_32_1
      & COMPUTE_OUTER_LOOP_stage_0_1 & (fsm_output[2]);
  assign and_152_rmff = COMPUTE_OUTER_LOOP_stage_0_6 & (~ CALC_SOFTMAX_LOOP_equal_tmp_20)
      & CALC_SOFTMAX_LOOP_equal_tmp_16 & (~ CALC_SOFTMAX_LOOP_equal_tmp_15) & CALC_SOFTMAX_LOOP_equal_tmp_14
      & (fsm_output[2]);
  assign and_163_rmff = CALC_SOFTMAX_LOOP_asn_itm & (~ exit_COMPUTE_OUTER_LOOP_sva_1)
      & COMPUTE_OUTER_LOOP_stage_0_1 & (fsm_output[3]);
  assign and_189_rmff = and_dcpl_87 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_0)
      & (~ CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_3) & (fsm_output[3]);
  assign COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_nor_cse = ~(or_dcpl_41 | (fsm_output[3]));
  assign or_78_nl = CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_3 | lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_0
      | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_1) | exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_3;
  assign mux_34_nl = MUX_s_1_2_2(not_tmp_75, or_dcpl_41, or_78_nl);
  assign COMPUTE_OUTER_LOOP_nor_2_seb = ~(and_191_cse | and_192_cse | mux_34_nl);
  assign and_210_rmff = and_dcpl_87 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_0)
      & CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_3 & (fsm_output[3]);
  assign or_82_nl = (~ CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_3) |
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_0 | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_1)
      | exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_3;
  assign mux_35_nl = MUX_s_1_2_2(not_tmp_75, or_dcpl_41, or_82_nl);
  assign COMPUTE_OUTER_LOOP_nor_1_seb = ~(and_191_cse | and_192_cse | mux_35_nl);
  assign COMPUTE_OUTER_LOOP_and_cse = compute_kernel_wen & (~((~ (fsm_output[2]))
      | (~ COMPUTE_OUTER_LOOP_stage_0_6) | CALC_SOFTMAX_LOOP_equal_tmp_20 | (~ CALC_SOFTMAX_LOOP_equal_tmp_16)
      | CALC_SOFTMAX_LOOP_equal_tmp_15 | (~ CALC_SOFTMAX_LOOP_equal_tmp_14)));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_and_cse = compute_kernel_wen
      & ((SUM_EXP_LOOP_acc_1_tmp!=74'b00000000000000000000000000000000000000000000000000000000000000000000000000))
      & and_dcpl_7 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_2_1) & CALC_SOFTMAX_LOOP_equal_tmp_10_2
      & (fsm_output[2]);
  assign CALC_SOFTMAX_LOOP_and_cse = compute_kernel_wen & (~((~((fsm_output[5]) |
      (fsm_output[2]))) | ((~ COMPUTE_OUTER_LOOP_stage_0_1) & (fsm_output[2]))));
  assign and_121_m1c = (COMPUTE_OUTER_LOOP_stage_0 | COMPUTE_OUTER_LOOP_stage_0_1)
      & (~ COMPUTE_OUTER_LOOP_asn_6_itm_2) & COMPUTE_OUTER_LOOP_stage_0_3;
  assign or_8_cse = (~ COMPUTE_OUTER_LOOP_stage_0_2) | COMPUTE_OUTER_LOOP_asn_6_itm_1;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_and_6_rgt
      = ((CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_itm & and_121_m1c) | (and_dcpl_108
      & COMPUTE_OUTER_LOOP_stage_0_3 & CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_itm))
      & (fsm_output[2]);
  assign COMPUTE_OUTER_LOOP_and_4_cse = compute_kernel_wen & (or_tmp_47 | (fsm_output[3]));
  assign CALC_SOFTMAX_LOOP_i_and_4_cse = compute_kernel_wen & (fsm_output[3]);
  assign or_173_tmp = or_dcpl_6 | (~(COMPUTE_OUTER_LOOP_stage_0_1 & (CALC_SOFTMAX_LOOP_acc_1_tmp[7])));
  assign CALC_SOFTMAX_LOOP_and_57_cse = compute_kernel_wen & ((~ CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_1)
      | (fsm_output[3]));
  assign CALC_SOFTMAX_LOOP_and_79_cse = compute_kernel_wen & (CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_1
      | (fsm_output[3]));
  assign CALC_SOFTMAX_LOOP_i_and_rgt = (~ CALC_SOFTMAX_LOOP_and_7_tmp) & and_138_m1c
      & (~ (fsm_output[3]));
  assign CALC_SOFTMAX_LOOP_i_and_1_rgt = CALC_SOFTMAX_LOOP_and_7_tmp & and_138_m1c
      & (~ (fsm_output[3]));
  assign and_140_rgt = or_dcpl_6 & (~((SUM_EXP_LOOP_acc_2_tmp[7]) & (CALC_EXP_LOOP_acc_1_tmp[7])))
      & COMPUTE_OUTER_LOOP_stage_0_1 & (~ (fsm_output[3]));
  assign CALC_SOFTMAX_LOOP_and_88_cse = compute_kernel_wen & (~ (fsm_output[3]));
  assign or_414_tmp = exit_COMPUTE_OUTER_LOOP_sva_1 | (~ CALC_SOFTMAX_LOOP_and_10_itm);
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_and_4_rgt
      = ~(or_414_tmp | (fsm_output[3]));
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_and_3_rgt
      = CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_itm & (~ or_162_tmp) & or_414_tmp
      & (~ (fsm_output[3]));
  assign and_615_rgt = or_162_tmp & or_414_tmp & (~ (fsm_output[3]));
  assign CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx1 = MUX_v_7_2_2(CALC_SOFTMAX_LOOP_i_7_0_lpi_2_dfm_2_6_0,
      CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0, or_8_cse);
  assign CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0 = MUX_v_5_2_2((CALC_SOFTMAX_LOOP_i_7_0_lpi_2_dfm_2_6_0[4:0]),
      (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[4:0]), or_8_cse);
  assign CALC_SOFTMAX_LOOP_equal_tmp_44_mx1w0 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b01011);
  assign CALC_SOFTMAX_LOOP_equal_tmp_40_mx1w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b00111);
  assign CALC_EXP_LOOP_and_svs_mx1w2 = (CALC_EXP_LOOP_acc_1_tmp[7]) & (SUM_EXP_LOOP_acc_2_tmp[7]);
  assign exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_1 = (~ COMPUTE_OUTER_LOOP_acc_itm_32_1)
      & exitL_exit_CALC_SOFTMAX_LOOP_sva;
  assign CALC_SOFTMAX_LOOP_equal_tmp_39_mx1w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[4:0]==5'b00110);
  assign CALC_SOFTMAX_LOOP_equal_tmp_57_mx1w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[4:0]==5'b11000);
  assign CALC_SOFTMAX_LOOP_equal_tmp_53_mx1w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[4:0]==5'b10100);
  assign CALC_SOFTMAX_LOOP_equal_tmp_51_mx1w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[4:0]==5'b10010);
  assign CALC_SOFTMAX_LOOP_equal_tmp_50_mx1w2 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[4:0]==5'b10001);
  assign CALC_SOFTMAX_LOOP_equal_tmp_49_mx1w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[4])
      & CALC_SOFTMAX_LOOP_nor_14_itm;
  assign CALC_SOFTMAX_LOOP_equal_tmp_45_mx1w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[4:0]==5'b01100);
  assign CALC_SOFTMAX_LOOP_equal_tmp_43_mx1w2 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[4:0]==5'b01010);
  assign CALC_SOFTMAX_LOOP_equal_tmp_42_mx1w2 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[4:0]==5'b01001);
  assign CALC_SOFTMAX_LOOP_equal_tmp_38_mx1w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[4:0]==5'b00101);
  assign CALC_SOFTMAX_LOOP_equal_tmp_37_mx1w0 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[2])
      & CALC_SOFTMAX_LOOP_nor_28_itm;
  assign CALC_SOFTMAX_LOOP_equal_tmp_36_mx1w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[4:0]==5'b00011);
  assign CALC_SOFTMAX_LOOP_equal_tmp_2_mx1w0 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[0])
      & CALC_SOFTMAX_LOOP_nor_25_itm;
  assign nl_COMPUTE_OUTER_LOOP_acc_nl = ({1'b1 , (~ COMPUTE_OUTER_LOOP_s_31_7_sva)
      , (~ (conf_info_crt_1_sva[6:0]))}) + 33'b000000000000000000000000000000001;
  assign COMPUTE_OUTER_LOOP_acc_nl = nl_COMPUTE_OUTER_LOOP_acc_nl[32:0];
  assign COMPUTE_OUTER_LOOP_acc_itm_32_1 = readslicef_33_1_32(COMPUTE_OUTER_LOOP_acc_nl);
  assign CALC_SOFTMAX_LOOP_equal_tmp_46_mx1w0 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b01101);
  assign CALC_SOFTMAX_LOOP_equal_tmp_47_mx1w0 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b01110);
  assign CALC_SOFTMAX_LOOP_equal_tmp_48_mx1w0 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b01111);
  assign CALC_SOFTMAX_LOOP_equal_tmp_52_mx1w0 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b10011);
  assign CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_6_0_mx1 = MUX_v_7_2_2(CALC_SOFTMAX_LOOP_i_7_0_lpi_2_dfm_2_6_0,
      (signext_7_1(~ COMPUTE_OUTER_LOOP_acc_itm_32_1)), exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign CALC_SOFTMAX_LOOP_nor_26_itm_mx1w0 = ~((CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0[4])
      | (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0[3]) | (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0[2])
      | (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0[0]));
  assign CALC_SOFTMAX_LOOP_nor_32_itm_mx1w1 = ~((CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0[4])
      | (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0[2]) | (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0[1])
      | (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0[0]));
  assign nl_SUM_EXP_LOOP_acc_1_tmp = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_2_dfm_1
      + conv_u2u_67_74(operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1);
  assign SUM_EXP_LOOP_acc_1_tmp = nl_SUM_EXP_LOOP_acc_1_tmp[73:0];
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = conv_u2u_19_19(({ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_itm_1
      , 1'b0 , ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_1_itm_1})
      * ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_32_14_11_0_1_itm_1);
  assign COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_and_4_mx0w0 = lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_1
      & (~ COMPUTE_OUTER_LOOP_acc_itm_32_1);
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_1_mx0 = MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_1,
      COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_and_4_mx0w0, exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_and_3_mx0w0 = lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_0
      & (~ COMPUTE_OUTER_LOOP_acc_itm_32_1);
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_0_mx0 = MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_0,
      COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_and_3_mx0w0, exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign nl_CALC_SOFTMAX_LOOP_acc_1_tmp = conv_u2u_7_8(CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx1)
      + 8'b00000001;
  assign CALC_SOFTMAX_LOOP_acc_1_tmp = nl_CALC_SOFTMAX_LOOP_acc_1_tmp[7:0];
  assign CALC_SOFTMAX_LOOP_equal_tmp_66 = lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_1_mx0
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_0_mx0);
  assign CALC_SOFTMAX_LOOP_or_tmp_1 = (lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_0_mx0
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_1_mx0)) | (~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_1_mx0
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_0_mx0));
  assign CALC_SOFTMAX_LOOP_equal_tmp_67 = lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_1_mx0
      & lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_0_mx0;
  assign CALC_SOFTMAX_LOOP_mux_183_nl = MUX_s_1_2_2((~ (CALC_SOFTMAX_LOOP_acc_1_tmp[7])),
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_1, CALC_SOFTMAX_LOOP_equal_tmp_67);
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_4_1_1 = (CALC_SOFTMAX_LOOP_mux_183_nl
      & (~ CALC_SOFTMAX_LOOP_and_4_ssc_1)) | CALC_SOFTMAX_LOOP_and_5_ssc_1;
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_4_0_1 = (lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_0_mx0
      & (~(CALC_SOFTMAX_LOOP_and_5_ssc_1 | CALC_SOFTMAX_LOOP_equal_tmp_66))) | CALC_SOFTMAX_LOOP_and_4_ssc_1;
  assign nl_CALC_EXP_LOOP_acc_1_tmp = conv_u2u_7_8(CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_6_0_mx1)
      + 8'b00000001;
  assign CALC_EXP_LOOP_acc_1_tmp = nl_CALC_EXP_LOOP_acc_1_tmp[7:0];
  assign CALC_SOFTMAX_LOOP_mux_184_nl = MUX_v_7_2_2(SUM_EXP_LOOP_i_7_0_lpi_2_6_0,
      (signext_7_1(~ COMPUTE_OUTER_LOOP_acc_itm_32_1)), exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign nl_SUM_EXP_LOOP_acc_2_tmp = conv_u2u_7_8(CALC_SOFTMAX_LOOP_mux_184_nl) +
      8'b00000001;
  assign SUM_EXP_LOOP_acc_2_tmp = nl_SUM_EXP_LOOP_acc_2_tmp[7:0];
  assign CALC_SOFTMAX_LOOP_and_4_ssc_1 = (~ CALC_EXP_LOOP_and_svs_mx1w2) & CALC_SOFTMAX_LOOP_or_tmp_1;
  assign CALC_SOFTMAX_LOOP_and_5_ssc_1 = CALC_EXP_LOOP_and_svs_mx1w2 & CALC_SOFTMAX_LOOP_or_tmp_1;
  assign CALC_SOFTMAX_LOOP_equal_tmp_64_mx0w0 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b11111);
  assign CALC_SOFTMAX_LOOP_equal_tmp_63_mx0w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b11110);
  assign CALC_SOFTMAX_LOOP_equal_tmp_62_mx0w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b11101);
  assign CALC_SOFTMAX_LOOP_equal_tmp_61_mx0w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b11100);
  assign CALC_SOFTMAX_LOOP_equal_tmp_60_mx0w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b11011);
  assign CALC_SOFTMAX_LOOP_equal_tmp_59_mx0w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b11010);
  assign CALC_SOFTMAX_LOOP_equal_tmp_58_mx0w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b11001);
  assign CALC_SOFTMAX_LOOP_equal_tmp_56_mx0w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b10111);
  assign CALC_SOFTMAX_LOOP_equal_tmp_55_mx0w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b10110);
  assign CALC_SOFTMAX_LOOP_equal_tmp_54_mx0w1 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0==5'b10101);
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_nl
      = MUX_v_8_8_2(8'b00011100, 8'b01001011, 8'b01101100, 8'b10000100, 8'b10010111,
      8'b10100110, 8'b10110011, 8'b10111100, ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_normalized_fixed_72_60_sva[12:10]);
  assign nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = $signed(({1'b1 , ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_nl}))
      * $signed(conv_u2s_10_11(ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_normalized_fixed_72_60_sva[9:0]));
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:0];
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_6_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[31:0]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[31:0]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_7_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[63:32]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[63:32]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_8_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[95:64]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[95:64]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_9_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[127:96]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[127:96]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_10_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[159:128]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[159:128]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_11_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[191:160]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[191:160]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_12_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[223:192]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[223:192]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_13_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[255:224]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[255:224]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_14_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[287:256]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[287:256]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_15_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[319:288]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[319:288]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_16_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[351:320]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[351:320]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_17_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[383:352]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[383:352]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_18_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[415:384]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[415:384]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_19_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[447:416]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[447:416]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_20_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[479:448]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[479:448]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_21_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[511:480]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[511:480]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_22_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[543:512]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[543:512]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_23_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[575:544]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[575:544]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_24_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[607:576]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[607:576]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_25_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[639:608]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[639:608]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_26_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[671:640]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[671:640]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_27_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[703:672]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[703:672]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_28_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[735:704]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[735:704]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_29_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[767:736]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[767:736]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_30_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[799:768]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[799:768]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_31_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[831:800]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[831:800]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_32_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[863:832]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[863:832]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_33_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[895:864]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[895:864]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_34_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[927:896]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[927:896]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_35_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[959:928]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[959:928]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_36_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[991:960]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[991:960]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_37_nl
      = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d[1023:992]),
      (COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d[1023:992]), CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[5]);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_5_nl
      = MUX_v_32_32_2(ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_6_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_7_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_8_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_9_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_10_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_11_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_12_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_13_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_14_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_15_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_16_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_17_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_18_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_19_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_20_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_21_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_22_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_23_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_24_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_25_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_26_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_27_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_28_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_29_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_30_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_31_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_32_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_33_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_34_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_35_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_36_nl,
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_37_nl,
      CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[4:0]);
  assign nl_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl
      = $signed(ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mux_5_nl)
      * $signed(16'b0101110001010101);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl
      = nl_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl[46:0];
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28
      = readslicef_47_19_28(ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl);
  assign CALC_SOFTMAX_LOOP_or_152 = CALC_SOFTMAX_LOOP_equal_tmp_2_3 | CALC_SOFTMAX_LOOP_equal_tmp_3_3
      | CALC_SOFTMAX_LOOP_equal_tmp_36_3 | CALC_SOFTMAX_LOOP_equal_tmp_37_2 | CALC_SOFTMAX_LOOP_equal_tmp_38_3
      | CALC_SOFTMAX_LOOP_equal_tmp_39_3 | CALC_SOFTMAX_LOOP_equal_tmp_40_3 | CALC_SOFTMAX_LOOP_equal_tmp_41_3
      | CALC_SOFTMAX_LOOP_equal_tmp_10_3 | CALC_SOFTMAX_LOOP_equal_tmp_11_3 | CALC_SOFTMAX_LOOP_equal_tmp_12_3
      | CALC_SOFTMAX_LOOP_equal_tmp_13_3 | CALC_SOFTMAX_LOOP_equal_tmp_14_3 | CALC_SOFTMAX_LOOP_equal_tmp_15_3
      | CALC_SOFTMAX_LOOP_equal_tmp_16_3 | CALC_SOFTMAX_LOOP_equal_tmp_17_3 | CALC_SOFTMAX_LOOP_equal_tmp_18_3
      | CALC_SOFTMAX_LOOP_equal_tmp_19_3 | CALC_SOFTMAX_LOOP_equal_tmp_20_3 | CALC_SOFTMAX_LOOP_equal_tmp_21_3
      | CALC_SOFTMAX_LOOP_equal_tmp_22_3 | CALC_SOFTMAX_LOOP_equal_tmp_23_3 | CALC_SOFTMAX_LOOP_equal_tmp_24_3
      | CALC_SOFTMAX_LOOP_equal_tmp_25_3 | CALC_SOFTMAX_LOOP_equal_tmp_26_3 | CALC_SOFTMAX_LOOP_equal_tmp_27_3
      | CALC_SOFTMAX_LOOP_equal_tmp_28_3 | CALC_SOFTMAX_LOOP_equal_tmp_29_3 | CALC_SOFTMAX_LOOP_equal_tmp_30_3
      | CALC_SOFTMAX_LOOP_equal_tmp_31_3 | CALC_SOFTMAX_LOOP_equal_tmp_32_3;
  assign or_dcpl_6 = exitL_exit_CALC_SOFTMAX_LOOP_sva | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_1);
  assign and_dcpl_7 = COMPUTE_OUTER_LOOP_stage_0_3 & (~ exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_2);
  assign and_dcpl_13 = COMPUTE_OUTER_LOOP_stage_0_2 & (~ COMPUTE_OUTER_LOOP_asn_6_itm_1);
  assign and_dcpl_87 = COMPUTE_OUTER_LOOP_stage_0_4 & (~ exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_3)
      & lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_1;
  assign or_dcpl_36 = (~ COMPUTE_OUTER_LOOP_stage_0_4) | exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_3
      | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_1);
  assign or_dcpl_41 = (~ COMPUTE_OUTER_LOOP_stage_0_5) | exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_4
      | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_4_1) | lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_4_0
      | (~ CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_4);
  assign not_tmp_75 = ~(COMPUTE_OUTER_LOOP_stage_0_4 | (~ or_dcpl_41));
  assign and_dcpl_108 = ~(COMPUTE_OUTER_LOOP_stage_0 | COMPUTE_OUTER_LOOP_stage_0_1);
  assign and_dcpl_113 = (~ exitL_exit_CALC_SOFTMAX_LOOP_sva) & lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_1;
  assign nor_13_nl = ~((~ (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_dfm_2_6_0[5])) | (~ COMPUTE_OUTER_LOOP_stage_0_2)
      | COMPUTE_OUTER_LOOP_asn_6_itm_1);
  assign or_168_nl = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_dfm_2_6_0[5]) | (~ COMPUTE_OUTER_LOOP_stage_0_2)
      | COMPUTE_OUTER_LOOP_asn_6_itm_1;
  assign mux_tmp_35 = MUX_s_1_2_2(nor_13_nl, or_168_nl, CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[5]);
  assign and_dcpl_114 = (~ mux_tmp_35) & and_dcpl_113;
  assign and_dcpl_115 = mux_tmp_35 & and_dcpl_113;
  assign and_dcpl_118 = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[5]) & CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm;
  assign or_tmp_47 = (fsm_output[1]) | (fsm_output[4]);
  assign and_191_cse = or_dcpl_41 & (fsm_output[3]);
  assign and_192_cse = ~((fsm_output[3:2]!=2'b00));
  assign and_239_cse = exitL_exit_CALC_SOFTMAX_LOOP_sva & (~ COMPUTE_OUTER_LOOP_acc_itm_32_1)
      & COMPUTE_OUTER_LOOP_stage_0_1 & (fsm_output[2]);
  assign COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_mux_7_rmff = CALC_SOFTMAX_LOOP_nor_1_itm
      & (~ (fsm_output[3]));
  assign CALC_SOFTMAX_LOOP_and_7_tmp = CALC_SOFTMAX_LOOP_equal_tmp_66 & (~ exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_1);
  assign and_138_m1c = (and_dcpl_113 | CALC_EXP_LOOP_and_svs_mx1w2) & COMPUTE_OUTER_LOOP_stage_0_1;
  assign or_162_tmp = COMPUTE_OUTER_LOOP_asn_6_itm_2 | (~ COMPUTE_OUTER_LOOP_stage_0_3);
  assign CALC_SOFTMAX_LOOP_mul_cmp_b = ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_2;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d
      = operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d
      = CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d
      = CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_6_0;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff
      = and_dcpl_7 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_2_1) & (fsm_output[2]);
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = and_dcpl_13 & lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_1 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_0)
      & (fsm_output[3]);
  assign COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_or_1_nl = (CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[6])
      | (fsm_output[3]);
  assign COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_adra_d = {(~ (fsm_output[3]))
      , COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_or_1_nl};
  assign COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_da_d = {(plm_in_cnsi_idat_mxwt[1023:0])
      , (plm_in_cnsi_idat_mxwt[3071:2048])};
  assign COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_wea_d = {{1{and_163_rmff}},
      and_163_rmff};
  assign and_166_nl = and_dcpl_13 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_1)
      & (~ CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_3_itm) & (fsm_output[2]);
  assign COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d
      = {1'b0 , and_166_nl};
  assign COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d
      = {{1{and_163_rmff}}, and_163_rmff};
  assign COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_and_nl = (CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0[6])
      & (~ (fsm_output[3]));
  assign COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_adra_d = {(fsm_output[3])
      , COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_and_nl};
  assign COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_da_d = {(plm_in_cnsi_idat_mxwt[4095:3072])
      , (plm_in_cnsi_idat_mxwt[2047:1024])};
  assign COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_wea_d = {{1{and_163_rmff}},
      and_163_rmff};
  assign and_178_nl = and_dcpl_13 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_1)
      & CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_3_itm & (fsm_output[2]);
  assign COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d
      = {1'b0 , and_178_nl};
  assign COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d
      = {{1{and_163_rmff}}, and_163_rmff};
  assign COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_or_5_cse = CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_3_itm_2
      | (~ (fsm_output[3]));
  assign COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_adra_d = {COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_or_5_cse
      , COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_mux_7_rmff};
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[1023:992]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_32_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_1_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[991:960]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_31_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_2_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[959:928]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_30_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_3_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[927:896]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_29_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_4_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[895:864]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_28_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_5_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[863:832]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_27_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_6_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[831:800]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_26_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_7_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[799:768]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_25_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_8_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[767:736]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_24_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_9_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[735:704]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_23_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_10_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[703:672]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_22_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_11_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[671:640]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_21_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_12_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[639:608]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_20_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_13_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[607:576]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_19_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_14_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[575:544]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_18_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_15_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[543:512]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_17_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_16_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[511:480]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_16_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_17_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[479:448]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_15_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_18_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[447:416]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_14_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_19_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[415:384]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_13_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_20_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[383:352]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_12_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_21_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[351:320]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_11_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_22_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[319:288]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_10_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_23_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[287:256]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_41_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_24_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[255:224]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_40_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_25_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[223:192]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_39_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_26_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[191:160]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_38_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_27_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[159:128]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_37_2);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_28_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[127:96]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_36_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_29_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[95:64]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_3_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_30_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[63:32]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_2_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_31_nl = MUX_v_32_2_2((CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]),
      (COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[31:0]), CALC_SOFTMAX_LOOP_or_152);
  assign COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_da_d = {CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_1_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_2_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_3_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_4_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_5_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_6_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_7_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_8_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_9_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_10_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_11_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_12_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_13_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_14_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_15_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_16_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_17_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_18_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_19_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_20_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_21_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_22_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_23_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_24_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_25_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_26_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_27_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_28_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_29_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_30_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_31_nl};
  assign COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_wea_d = {and_189_rmff ,
      1'b0};
  assign COMPUTE_OUTER_LOOP_and_9_nl = COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_nor_cse
      & COMPUTE_OUTER_LOOP_nor_2_seb;
  assign COMPUTE_OUTER_LOOP_and_13_nl = (~((or_dcpl_36 | lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_0
      | CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_3) & (~ or_dcpl_41)
      & (fsm_output[2]))) & COMPUTE_OUTER_LOOP_nor_2_seb;
  assign COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d
      = {COMPUTE_OUTER_LOOP_and_9_nl , COMPUTE_OUTER_LOOP_and_13_nl};
  assign COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d
      = {and_189_rmff , 1'b0};
  assign COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_adra_d = {COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_or_5_cse
      , COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_mux_7_rmff};
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_32_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[1023:992]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_32_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_33_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[991:960]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_31_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_34_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[959:928]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_30_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_35_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[927:896]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_29_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_36_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[895:864]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_28_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_37_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[863:832]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_27_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_38_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[831:800]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_26_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_39_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[799:768]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_25_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_40_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[767:736]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_24_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_41_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[735:704]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_23_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_42_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[703:672]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_22_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_43_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[671:640]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_21_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_44_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[639:608]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_20_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_45_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[607:576]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_19_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_46_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[575:544]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_18_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_47_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[543:512]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_17_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_48_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[511:480]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_16_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_49_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[479:448]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_15_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_50_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[447:416]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_14_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_51_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[415:384]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_13_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_52_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[383:352]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_12_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_53_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[351:320]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_11_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_54_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[319:288]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_10_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_55_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[287:256]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_41_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_56_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[255:224]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_40_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_57_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[223:192]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_39_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_58_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[191:160]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_38_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_59_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[159:128]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_37_2);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_60_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[127:96]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_36_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_61_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[95:64]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_3_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_62_nl = MUX_v_32_2_2((COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[63:32]),
      (CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]), CALC_SOFTMAX_LOOP_equal_tmp_2_3);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_63_nl = MUX_v_32_2_2((CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]),
      (COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[31:0]), CALC_SOFTMAX_LOOP_or_152);
  assign COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_da_d = {CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_32_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_33_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_34_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_35_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_36_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_37_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_38_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_39_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_40_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_41_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_42_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_43_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_44_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_45_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_46_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_47_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_48_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_49_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_50_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_51_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_52_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_53_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_54_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_55_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_56_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_57_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_58_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_59_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_60_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_61_nl , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_62_nl
      , CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_63_nl};
  assign COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_wea_d = {and_210_rmff ,
      1'b0};
  assign COMPUTE_OUTER_LOOP_and_10_nl = COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_nor_cse
      & COMPUTE_OUTER_LOOP_nor_1_seb;
  assign COMPUTE_OUTER_LOOP_and_14_nl = (~((or_dcpl_36 | lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_0
      | (~ CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_3)) & (~ or_dcpl_41)
      & (fsm_output[2]))) & COMPUTE_OUTER_LOOP_nor_1_seb;
  assign COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d
      = {COMPUTE_OUTER_LOOP_and_10_nl , COMPUTE_OUTER_LOOP_and_14_nl};
  assign COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d
      = {and_210_rmff , 1'b0};
  always @(posedge clk) begin
    if ( compute_kernel_wen ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_2
          <= MUX_v_94_2_2(ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_2,
          ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_or_nl,
          and_247_nl);
      tmp_4_sva_1 <= COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[2047:1024];
      tmp_3_sva_1 <= COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[2047:1024];
      ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_2_itm_1
          <= MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28[11:10]);
      ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_3_itm_1
          <= MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28[11:10]);
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_32_14_18_12_itm_1
          <= ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28[18:12];
      ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_itm_1
          <= MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28[11:10]);
      ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_1_itm_1
          <= MUX_v_3_4_2(3'b010, 3'b110, 3'b001, 3'b101, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28[11:10]);
      ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_slc_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_input_inter_32_14_11_0_1_itm_1
          <= ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28[9:0];
      COMPUTE_OUTER_LOOP_s_31_7_sva <= MUX1HOT_v_25_4_2((conf_info_crt_1_sva[31:7]),
          (conf_info[31:7]), (z_out_1[24:0]), COMPUTE_OUTER_LOOP_s_31_7_sva, {COMPUTE_OUTER_LOOP_s_and_nl
          , (fsm_output[1]) , COMPUTE_OUTER_LOOP_s_and_2_nl , COMPUTE_OUTER_LOOP_s_or_nl});
      conf_info_crt_1_sva <= MUX_v_64_2_2(conf_info, conf_info_crt_1_sva, or_269_nl);
      CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_3_itm_2 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_3_itm_2,
          CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_3_itm_1, fsm_output[3]);
      COMPUTE_BATCH_LOOP_b_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          COMPUTE_BATCH_LOOP_b_mux_nl, softmax_softmax_not_nl);
      CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_5_itm <= CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[6];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_input_ready_channel_Push_mioi_oswt_cse <= 1'b0;
      reg_output_ready_channel_Pop_mioi_oswt_cse <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm <= 1'b0;
      exitL_exit_CALC_SOFTMAX_LOOP_sva <= 1'b0;
      CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_3 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_0 <= 1'b0;
      exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_3 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_2_1 <= 1'b0;
      exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_2 <= 1'b0;
      CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0 <= 7'b0000000;
      CALC_SOFTMAX_LOOP_asn_itm_1 <= 1'b0;
      COMPUTE_OUTER_LOOP_stage_0 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_32_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_31_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_30_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_29_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_28_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_27_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_26_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_25_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_24_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_23_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_22_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_21_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_20_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_19_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_18_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_17_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_16_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_15_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_14_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_13_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_12_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_11_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_10_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_3_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_2_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_41_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_40_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_39_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_38_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_37_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_36_3 <= 1'b0;
      COMPUTE_OUTER_LOOP_stage_0_6 <= 1'b0;
      exit_COMPUTE_OUTER_LOOP_sva_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_itm <= 1'b0;
      CALC_SOFTMAX_LOOP_and_10_itm <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_14 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_15 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_16 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_20 <= 1'b0;
      CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_6_0 <= 7'b0000000;
      CALC_SOFTMAX_LOOP_nor_1_itm <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_0 <= 1'b0;
      CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_3_itm <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_32 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_31 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_30 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_29 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_28 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_27 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_26 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_24 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_23 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_22 <= 1'b0;
      CALC_SOFTMAX_LOOP_nor_14_itm <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_64 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm <= 1'b0;
    end
    else if ( compute_kernel_wen ) begin
      reg_input_ready_channel_Push_mioi_oswt_cse <= and_150_rmff;
      reg_output_ready_channel_Pop_mioi_oswt_cse <= and_152_rmff;
      CALC_SOFTMAX_LOOP_asn_itm <= COMPUTE_OUTER_LOOP_mux_33_nl | or_tmp_47;
      exitL_exit_CALC_SOFTMAX_LOOP_sva <= COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_mux_nl
          | or_tmp_47;
      CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_3,
          CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2, fsm_output[3]);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_1,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_2_1, fsm_output[3]);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_0 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_0,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_2_0, fsm_output[3]);
      exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_3 <= MUX_s_1_2_2(exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_3,
          exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_2, fsm_output[3]);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_2_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_2_1,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_1, fsm_output[3]);
      exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_2 <= MUX_s_1_2_2(exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_2,
          COMPUTE_OUTER_LOOP_asn_6_itm_1, fsm_output[3]);
      CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0 <= MUX1HOT_v_7_3_2(CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0,
          CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0, CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_6_0,
          {CALC_EXP_LOOP_i_CALC_EXP_LOOP_i_nor_nl , CALC_EXP_LOOP_i_and_1_nl , (fsm_output[3])});
      CALC_SOFTMAX_LOOP_asn_itm_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_mux1h_22_nl, CALC_SOFTMAX_LOOP_asn_itm,
          fsm_output[3]);
      COMPUTE_OUTER_LOOP_stage_0 <= (COMPUTE_OUTER_LOOP_stage_0 | (~((fsm_output[3])
          | ((COMPUTE_OUTER_LOOP_acc_itm_32_1 | (~ exitL_exit_CALC_SOFTMAX_LOOP_sva)
          | (~ COMPUTE_OUTER_LOOP_stage_0_1)) & (fsm_output[2]))))) & (~((fsm_output[0])
          | (fsm_output[5]) | and_239_cse));
      CALC_SOFTMAX_LOOP_equal_tmp_32_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_32_3,
          CALC_SOFTMAX_LOOP_mux_14_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_31_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_31_3,
          CALC_SOFTMAX_LOOP_mux_16_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_30_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_30_3,
          CALC_SOFTMAX_LOOP_mux_18_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_29_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_29_3,
          CALC_SOFTMAX_LOOP_mux_20_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_28_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_28_3,
          CALC_SOFTMAX_LOOP_mux_22_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_27_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_27_3,
          CALC_SOFTMAX_LOOP_mux_24_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_26_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_26_3,
          CALC_SOFTMAX_LOOP_mux_26_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_25_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_25_3,
          CALC_SOFTMAX_LOOP_mux_28_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_24_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_24_3,
          CALC_SOFTMAX_LOOP_mux_30_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_23_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_23_3,
          CALC_SOFTMAX_LOOP_mux_32_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_22_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_22_3,
          CALC_SOFTMAX_LOOP_mux_34_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_21_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_21_3,
          CALC_SOFTMAX_LOOP_mux_36_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_20_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_20_3,
          CALC_SOFTMAX_LOOP_mux_38_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_19_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_19_3,
          CALC_SOFTMAX_LOOP_mux_40_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_18_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_18_3,
          CALC_SOFTMAX_LOOP_mux_42_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_17_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_17_3,
          CALC_SOFTMAX_LOOP_mux_44_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_16_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_16_3,
          CALC_SOFTMAX_LOOP_mux_46_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_15_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_15_3,
          CALC_SOFTMAX_LOOP_mux_48_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_14_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_14_3,
          CALC_SOFTMAX_LOOP_mux_50_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_13_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_13_3,
          CALC_SOFTMAX_LOOP_mux_52_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_12_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_12_3,
          CALC_SOFTMAX_LOOP_mux_54_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_11_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_11_3,
          CALC_SOFTMAX_LOOP_mux_56_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_10_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_10_3,
          CALC_SOFTMAX_LOOP_mux_58_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_3_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_3_3,
          CALC_SOFTMAX_LOOP_mux_60_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_2_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_2_3,
          CALC_SOFTMAX_LOOP_mux_62_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_41_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_41_3,
          CALC_SOFTMAX_LOOP_mux_64_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_40_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_40_3,
          CALC_SOFTMAX_LOOP_mux_66_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_39_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_39_3,
          CALC_SOFTMAX_LOOP_mux_68_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_38_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_38_3,
          CALC_SOFTMAX_LOOP_mux_70_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_37_2 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_37_2,
          CALC_SOFTMAX_LOOP_mux_72_nl, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_36_3 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_36_3,
          CALC_SOFTMAX_LOOP_mux_74_nl, fsm_output[3]);
      COMPUTE_OUTER_LOOP_stage_0_6 <= COMPUTE_OUTER_LOOP_mux_32_nl & (~ or_tmp_47);
      exit_COMPUTE_OUTER_LOOP_sva_1 <= MUX_s_1_2_2((~ COMPUTE_OUTER_LOOP_acc_itm_32_1),
          exit_COMPUTE_OUTER_LOOP_sva_1, fsm_output[3]);
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_itm <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_nl,
          CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_itm_1, fsm_output[3]);
      CALC_SOFTMAX_LOOP_and_10_itm <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_and_10_nl, CALC_SOFTMAX_LOOP_asn_3_itm,
          fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_14 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_mux_164_nl,
          CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_4, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_15 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_mux_166_nl,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_4_0, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_16 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_mux_168_nl,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_4_1, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_20 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_mux_170_nl,
          exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_4, fsm_output[3]);
      CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_6_0 <= MUX_v_7_2_2(CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_6_0_mx1,
          CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_1_6_0, fsm_output[3]);
      CALC_SOFTMAX_LOOP_nor_1_itm <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_mux1h_228_nl,
          CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_3_itm_1, fsm_output[3]);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_1_mx0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_0_mx0;
      CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm <= CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx1[5];
      CALC_SOFTMAX_LOOP_asn_3_itm <= exitL_exit_CALC_SOFTMAX_LOOP_sva;
      CALC_SOFTMAX_LOOP_equal_tmp_32 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_64_mx0w0,
          CALC_SOFTMAX_LOOP_equal_tmp_63_mx0w1, mux_tmp_35);
      CALC_SOFTMAX_LOOP_equal_tmp_31 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_63_mx0w1,
          CALC_SOFTMAX_LOOP_equal_tmp_62_mx0w1, mux_tmp_35);
      CALC_SOFTMAX_LOOP_equal_tmp_30 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_62_mx0w1,
          CALC_SOFTMAX_LOOP_equal_tmp_61_mx0w1, mux_tmp_35);
      CALC_SOFTMAX_LOOP_equal_tmp_29 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_61_mx0w1,
          CALC_SOFTMAX_LOOP_equal_tmp_60_mx0w1, mux_tmp_35);
      CALC_SOFTMAX_LOOP_equal_tmp_28 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_60_mx0w1,
          CALC_SOFTMAX_LOOP_equal_tmp_59_mx0w1, mux_tmp_35);
      CALC_SOFTMAX_LOOP_equal_tmp_27 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_59_mx0w1,
          CALC_SOFTMAX_LOOP_equal_tmp_58_mx0w1, mux_tmp_35);
      CALC_SOFTMAX_LOOP_equal_tmp_26 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_58_mx0w1,
          CALC_SOFTMAX_LOOP_equal_tmp_56_mx0w1, mux_tmp_35);
      CALC_SOFTMAX_LOOP_equal_tmp_24 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_56_mx0w1,
          CALC_SOFTMAX_LOOP_equal_tmp_55_mx0w1, mux_tmp_35);
      CALC_SOFTMAX_LOOP_equal_tmp_23 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_55_mx0w1,
          CALC_SOFTMAX_LOOP_equal_tmp_54_mx0w1, mux_tmp_35);
      CALC_SOFTMAX_LOOP_equal_tmp_22 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_54_mx0w1,
          CALC_SOFTMAX_LOOP_equal_tmp_52_mx1w0, mux_tmp_35);
      CALC_SOFTMAX_LOOP_nor_14_itm <= ~((CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0[3:0]!=4'b0000));
      CALC_SOFTMAX_LOOP_equal_tmp_64 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_40_mx1w1,
          CALC_SOFTMAX_LOOP_equal_tmp_64_mx0w0, mux_tmp_35);
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm <= CALC_SOFTMAX_LOOP_acc_1_tmp[7];
    end
  end
  always @(posedge clk) begin
    if ( COMPUTE_OUTER_LOOP_and_cse ) begin
      plm_out_cnsi_idat_2047_1024 <= COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d[1023:0];
      plm_out_cnsi_idat_3071_2048 <= tmp_3_sva_1;
      plm_out_cnsi_idat_1023_0 <= COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d[1023:0];
      plm_out_cnsi_idat_4095_3072 <= tmp_4_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_and_cse ) begin
      ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm <= nl_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm[7:0];
      ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_normalized_fixed_72_60_sva
          <= operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm[72:60];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_0 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_1 <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_cse ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_0 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_4_0_1,
          COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_and_3_mx0w0, and_239_cse);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_4_1_1,
          COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_and_4_mx0w0, and_239_cse);
    end
  end
  always @(posedge clk) begin
    if ( compute_kernel_wen & (((((~ CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_itm)
        & and_121_m1c) | (and_dcpl_108 & COMPUTE_OUTER_LOOP_stage_0_3 & (~ CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_itm)))
        & (fsm_output[2])) | ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_and_6_rgt)
        ) begin
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_2
          <= MUX_v_74_2_2(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_2_dfm_1,
          SUM_EXP_LOOP_acc_1_tmp, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_and_6_rgt);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      COMPUTE_OUTER_LOOP_stage_0_1 <= 1'b0;
      COMPUTE_OUTER_LOOP_stage_0_2 <= 1'b0;
      COMPUTE_OUTER_LOOP_stage_0_3 <= 1'b0;
      COMPUTE_OUTER_LOOP_stage_0_4 <= 1'b0;
      COMPUTE_OUTER_LOOP_stage_0_5 <= 1'b0;
    end
    else if ( COMPUTE_OUTER_LOOP_and_4_cse ) begin
      COMPUTE_OUTER_LOOP_stage_0_1 <= COMPUTE_OUTER_LOOP_stage_0 | (~ (fsm_output[3]));
      COMPUTE_OUTER_LOOP_stage_0_2 <= COMPUTE_OUTER_LOOP_stage_0_1 & (fsm_output[3]);
      COMPUTE_OUTER_LOOP_stage_0_3 <= COMPUTE_OUTER_LOOP_stage_0_2 & (fsm_output[3]);
      COMPUTE_OUTER_LOOP_stage_0_4 <= COMPUTE_OUTER_LOOP_stage_0_3 & (fsm_output[3]);
      COMPUTE_OUTER_LOOP_stage_0_5 <= COMPUTE_OUTER_LOOP_stage_0_4 & (fsm_output[3]);
    end
  end
  always @(posedge clk) begin
    if ( CALC_SOFTMAX_LOOP_i_and_4_cse ) begin
      CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_3_itm_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_5_itm,
          CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_3_itm, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_4 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_4_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_4_0 <= 1'b0;
      exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_4 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_2_0 <= 1'b0;
      COMPUTE_OUTER_LOOP_asn_6_itm_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_0 <= 1'b0;
      COMPUTE_OUTER_LOOP_asn_6_itm_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_and_10_itm_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_64_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_63_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_62_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_32_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_31_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_30_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_29_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_28_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_27_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_26_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_25_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_24_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_23_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_22_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_21_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_20_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_19_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_18_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_17_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_16_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_15_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_14_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_13_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_12_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_10_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_6_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_5_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_4_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_3_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_2_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_itm_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_and_10_itm_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_63_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_62_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_32_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_31_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_30_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_29_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_28_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_27_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_26_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_25_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_24_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_23_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_22_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_21_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_20_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_19_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_18_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_17_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_16_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_15_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_14_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_12_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_6_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_4_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_3_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_2_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_1 <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_i_and_4_cse ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_4 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_3;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_4_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_4_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_3_0;
      exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_4 <= exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_st_3;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_2_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_0;
      COMPUTE_OUTER_LOOP_asn_6_itm_2 <= COMPUTE_OUTER_LOOP_asn_6_itm_1;
      CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_1 <= CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_0;
      COMPUTE_OUTER_LOOP_asn_6_itm_1 <= COMPUTE_OUTER_LOOP_stage_0_6;
      CALC_SOFTMAX_LOOP_and_10_itm_2 <= CALC_SOFTMAX_LOOP_and_10_itm_1;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_3 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_2;
      CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2 <= CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_1;
      CALC_SOFTMAX_LOOP_equal_tmp_64_2 <= CALC_SOFTMAX_LOOP_equal_tmp_64_1;
      CALC_SOFTMAX_LOOP_equal_tmp_63_2 <= CALC_SOFTMAX_LOOP_equal_tmp_63_1;
      CALC_SOFTMAX_LOOP_equal_tmp_62_2 <= CALC_SOFTMAX_LOOP_equal_tmp_62_1;
      CALC_SOFTMAX_LOOP_equal_tmp_32_2 <= CALC_SOFTMAX_LOOP_equal_tmp_32_1;
      CALC_SOFTMAX_LOOP_equal_tmp_31_2 <= CALC_SOFTMAX_LOOP_equal_tmp_31_1;
      CALC_SOFTMAX_LOOP_equal_tmp_30_2 <= CALC_SOFTMAX_LOOP_equal_tmp_30_1;
      CALC_SOFTMAX_LOOP_equal_tmp_29_2 <= CALC_SOFTMAX_LOOP_equal_tmp_29_1;
      CALC_SOFTMAX_LOOP_equal_tmp_28_2 <= CALC_SOFTMAX_LOOP_equal_tmp_28_1;
      CALC_SOFTMAX_LOOP_equal_tmp_27_2 <= CALC_SOFTMAX_LOOP_equal_tmp_27_1;
      CALC_SOFTMAX_LOOP_equal_tmp_26_2 <= CALC_SOFTMAX_LOOP_equal_tmp_26_1;
      CALC_SOFTMAX_LOOP_equal_tmp_25_2 <= CALC_SOFTMAX_LOOP_equal_tmp_25_1;
      CALC_SOFTMAX_LOOP_equal_tmp_24_2 <= CALC_SOFTMAX_LOOP_equal_tmp_24_1;
      CALC_SOFTMAX_LOOP_equal_tmp_23_2 <= CALC_SOFTMAX_LOOP_equal_tmp_23_1;
      CALC_SOFTMAX_LOOP_equal_tmp_22_2 <= CALC_SOFTMAX_LOOP_equal_tmp_22_1;
      CALC_SOFTMAX_LOOP_equal_tmp_21_2 <= CALC_SOFTMAX_LOOP_equal_tmp_21_1;
      CALC_SOFTMAX_LOOP_equal_tmp_20_2 <= CALC_SOFTMAX_LOOP_equal_tmp_20_1;
      CALC_SOFTMAX_LOOP_equal_tmp_19_2 <= CALC_SOFTMAX_LOOP_equal_tmp_19_1;
      CALC_SOFTMAX_LOOP_equal_tmp_18_2 <= CALC_SOFTMAX_LOOP_equal_tmp_18_1;
      CALC_SOFTMAX_LOOP_equal_tmp_17_2 <= CALC_SOFTMAX_LOOP_equal_tmp_17_1;
      CALC_SOFTMAX_LOOP_equal_tmp_16_2 <= CALC_SOFTMAX_LOOP_equal_tmp_16_1;
      CALC_SOFTMAX_LOOP_equal_tmp_15_2 <= CALC_SOFTMAX_LOOP_equal_tmp_15_1;
      CALC_SOFTMAX_LOOP_equal_tmp_14_2 <= CALC_SOFTMAX_LOOP_equal_tmp_14_1;
      CALC_SOFTMAX_LOOP_equal_tmp_13_2 <= CALC_SOFTMAX_LOOP_equal_tmp_13_1;
      CALC_SOFTMAX_LOOP_equal_tmp_12_2 <= CALC_SOFTMAX_LOOP_equal_tmp_12_1;
      CALC_SOFTMAX_LOOP_equal_tmp_10_2 <= CALC_SOFTMAX_LOOP_equal_tmp_10_1;
      CALC_SOFTMAX_LOOP_equal_tmp_6_2 <= CALC_SOFTMAX_LOOP_equal_tmp_6_1;
      CALC_SOFTMAX_LOOP_equal_tmp_5_1 <= CALC_SOFTMAX_LOOP_equal_tmp_5;
      CALC_SOFTMAX_LOOP_equal_tmp_4_2 <= CALC_SOFTMAX_LOOP_equal_tmp_4_1;
      CALC_SOFTMAX_LOOP_equal_tmp_3_2 <= CALC_SOFTMAX_LOOP_equal_tmp_3_1;
      CALC_SOFTMAX_LOOP_equal_tmp_2_2 <= CALC_SOFTMAX_LOOP_equal_tmp_2_1;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_itm_1 <= CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_itm;
      CALC_SOFTMAX_LOOP_and_10_itm_1 <= CALC_SOFTMAX_LOOP_and_10_itm;
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_2 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_1;
      CALC_SOFTMAX_LOOP_equal_tmp_63_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_64,
          CALC_SOFTMAX_LOOP_equal_tmp_32, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm);
      CALC_SOFTMAX_LOOP_equal_tmp_62_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_31,
          CALC_SOFTMAX_LOOP_equal_tmp_39_mx1w1, nor_nl);
      CALC_SOFTMAX_LOOP_equal_tmp_32_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_32,
          CALC_SOFTMAX_LOOP_equal_tmp_27, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm);
      CALC_SOFTMAX_LOOP_equal_tmp_31_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_31,
          CALC_SOFTMAX_LOOP_equal_tmp_57_mx1w1, and_dcpl_118);
      CALC_SOFTMAX_LOOP_equal_tmp_30_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_30,
          CALC_SOFTMAX_LOOP_equal_tmp_26, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm);
      CALC_SOFTMAX_LOOP_equal_tmp_29_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_29,
          CALC_SOFTMAX_LOOP_equal_tmp_23, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm);
      CALC_SOFTMAX_LOOP_equal_tmp_28_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_28,
          CALC_SOFTMAX_LOOP_equal_tmp_53_mx1w1, and_dcpl_118);
      CALC_SOFTMAX_LOOP_equal_tmp_27_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_27,
          CALC_SOFTMAX_LOOP_equal_tmp_22, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm);
      CALC_SOFTMAX_LOOP_equal_tmp_26_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_26,
          CALC_SOFTMAX_LOOP_equal_tmp_51_mx1w1, and_dcpl_118);
      CALC_SOFTMAX_LOOP_equal_tmp_25_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_57_mx1w1,
          CALC_SOFTMAX_LOOP_equal_tmp_50_mx1w2, and_dcpl_118);
      CALC_SOFTMAX_LOOP_equal_tmp_24_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_24,
          CALC_SOFTMAX_LOOP_equal_tmp_49_mx1w1, and_dcpl_118);
      CALC_SOFTMAX_LOOP_equal_tmp_23_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_23,
          CALC_SOFTMAX_LOOP_equal_tmp_20, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm);
      CALC_SOFTMAX_LOOP_equal_tmp_22_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_22,
          CALC_SOFTMAX_LOOP_equal_tmp_16, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm);
      CALC_SOFTMAX_LOOP_equal_tmp_21_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_53_mx1w1,
          CALC_SOFTMAX_LOOP_equal_tmp_15, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm);
      CALC_SOFTMAX_LOOP_equal_tmp_20_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_20,
          CALC_SOFTMAX_LOOP_equal_tmp_45_mx1w1, and_dcpl_118);
      CALC_SOFTMAX_LOOP_equal_tmp_19_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_51_mx1w1,
          CALC_SOFTMAX_LOOP_equal_tmp_43_mx1w2, and_dcpl_118);
      CALC_SOFTMAX_LOOP_equal_tmp_18_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_50_mx1w2,
          CALC_SOFTMAX_LOOP_equal_tmp_42_mx1w2, and_dcpl_118);
      CALC_SOFTMAX_LOOP_equal_tmp_17_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_49_mx1w1,
          CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_41_nl, and_dcpl_118);
      CALC_SOFTMAX_LOOP_equal_tmp_16_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_16,
          CALC_SOFTMAX_LOOP_asn_itm_1, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm);
      CALC_SOFTMAX_LOOP_equal_tmp_15_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_15,
          CALC_SOFTMAX_LOOP_equal_tmp_39_mx1w1, and_dcpl_118);
      CALC_SOFTMAX_LOOP_equal_tmp_14_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_14,
          CALC_SOFTMAX_LOOP_equal_tmp_38_mx1w1, and_dcpl_118);
      CALC_SOFTMAX_LOOP_equal_tmp_12_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_asn_itm_1,
          CALC_SOFTMAX_LOOP_equal_tmp_36_mx1w1, and_dcpl_118);
      CALC_SOFTMAX_LOOP_equal_tmp_6_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_38_mx1w1,
          CALC_SOFTMAX_LOOP_equal_tmp_30, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm);
      CALC_SOFTMAX_LOOP_equal_tmp_4_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_36_mx1w1,
          CALC_SOFTMAX_LOOP_equal_tmp_28, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm);
      CALC_SOFTMAX_LOOP_equal_tmp_3_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_4_nl,
          CALC_SOFTMAX_LOOP_equal_tmp_24, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm);
      CALC_SOFTMAX_LOOP_equal_tmp_2_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_2_mx1w0,
          CALC_SOFTMAX_LOOP_equal_tmp_14, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm);
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm_1 <= CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_7_itm;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0 <= 7'b0000000;
    end
    else if ( compute_kernel_wen & (~(or_8_cse | (fsm_output[3]))) ) begin
      CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0 <= CALC_SOFTMAX_LOOP_i_7_0_lpi_2_dfm_2_6_0;
    end
  end
  always @(posedge clk) begin
    if ( compute_kernel_wen & COMPUTE_OUTER_LOOP_stage_0_1 & (~ (fsm_output[3]))
        ) begin
      SUM_EXP_LOOP_i_7_0_lpi_2_6_0 <= SUM_EXP_LOOP_acc_2_tmp[6:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_equal_tmp_11_2 <= 1'b0;
    end
    else if ( compute_kernel_wen & ((~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_2_1)
        | (fsm_output[3])) ) begin
      CALC_SOFTMAX_LOOP_equal_tmp_11_2 <= MUX_s_1_2_2(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_nl,
          CALC_SOFTMAX_LOOP_equal_tmp_11_1, fsm_output[3]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_equal_tmp_64_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_5 <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_57_cse ) begin
      CALC_SOFTMAX_LOOP_equal_tmp_64_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_10_nl,
          CALC_SOFTMAX_LOOP_equal_tmp_64, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_5 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_37_mx1w0,
          CALC_SOFTMAX_LOOP_equal_tmp_29, fsm_output[3]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_equal_tmp_13_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_equal_tmp_11_1 <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_79_cse ) begin
      CALC_SOFTMAX_LOOP_equal_tmp_13_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_37_mx1w0,
          CALC_SOFTMAX_LOOP_equal_tmp_45_mx1w1, fsm_output[3]);
      CALC_SOFTMAX_LOOP_equal_tmp_11_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_35_nl,
          CALC_SOFTMAX_LOOP_equal_tmp_43_mx1w2, fsm_output[3]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_equal_tmp_10_1 <= 1'b0;
    end
    else if ( compute_kernel_wen & ((lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_1
        & CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_1) | (fsm_output[3]))
        ) begin
      CALC_SOFTMAX_LOOP_equal_tmp_10_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_2_mx1w0,
          CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_68_nl, fsm_output[3]);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_i_7_0_lpi_2_dfm_2_6_0 <= 7'b0000000;
    end
    else if ( compute_kernel_wen & (CALC_SOFTMAX_LOOP_i_and_rgt | CALC_SOFTMAX_LOOP_i_and_1_rgt
        | and_140_rgt) ) begin
      CALC_SOFTMAX_LOOP_i_7_0_lpi_2_dfm_2_6_0 <= MUX1HOT_v_7_3_2((signext_7_1(~ CALC_EXP_LOOP_and_svs_mx1w2)),
          (CALC_SOFTMAX_LOOP_acc_1_tmp[6:0]), (CALC_EXP_LOOP_acc_1_tmp[6:0]), {CALC_SOFTMAX_LOOP_i_and_rgt
          , CALC_SOFTMAX_LOOP_i_and_1_rgt , and_140_rgt});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_nor_25_itm <= 1'b0;
      CALC_SOFTMAX_LOOP_nor_26_itm <= 1'b0;
      CALC_SOFTMAX_LOOP_nor_28_itm <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_88_cse ) begin
      CALC_SOFTMAX_LOOP_nor_25_itm <= ~((CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0[4:1]!=4'b0000));
      CALC_SOFTMAX_LOOP_nor_26_itm <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_nor_32_itm_mx1w1,
          CALC_SOFTMAX_LOOP_nor_26_itm_mx1w0, mux_tmp_35);
      CALC_SOFTMAX_LOOP_nor_28_itm <= ~((CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0[4])
          | (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0[3]) | (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0[1])
          | (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0_mx2_4_0[0]));
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_3_itm <= 1'b0;
    end
    else if ( compute_kernel_wen & (lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_1
        | (fsm_output[3])) ) begin
      CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_3_itm <= MUX_s_1_2_2((CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[6]),
          CALC_SOFTMAX_LOOP_nor_1_itm, fsm_output[3]);
    end
  end
  always @(posedge clk) begin
    if ( compute_kernel_wen & (ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_and_4_rgt
        | ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_and_3_rgt
        | and_615_rgt) ) begin
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_2_dfm_1
          <= MUX1HOT_v_74_3_2(({{73{exit_COMPUTE_OUTER_LOOP_sva_1}}, exit_COMPUTE_OUTER_LOOP_sva_1}),
          SUM_EXP_LOOP_acc_1_tmp, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_2,
          {ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_and_4_rgt
          , ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_and_3_rgt
          , and_615_rgt});
    end
  end
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_or_nl
      = MUX_v_94_2_2(operator_94_21_false_AC_TRN_AC_WRAP_rshift_itm, 94'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
      CALC_SOFTMAX_LOOP_equal_tmp_11_2);
  assign and_247_nl = (~((COMPUTE_OUTER_LOOP_stage_0 | COMPUTE_OUTER_LOOP_stage_0_2
      | COMPUTE_OUTER_LOOP_stage_0_1) & COMPUTE_OUTER_LOOP_asn_6_itm_2)) & COMPUTE_OUTER_LOOP_stage_0_3
      & CALC_SOFTMAX_LOOP_and_10_itm_2 & (fsm_output[3]);
  assign COMPUTE_OUTER_LOOP_mux_33_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_asn_itm, exitL_exit_CALC_SOFTMAX_LOOP_sva,
      fsm_output[3]);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_nl = ~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_4_1_1
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_4_0_1);
  assign COMPUTE_OUTER_LOOP_and_16_nl = COMPUTE_OUTER_LOOP_stage_0_1 & (fsm_output[2]);
  assign COMPUTE_OUTER_LOOP_COMPUTE_OUTER_LOOP_mux_nl = MUX_s_1_2_2(exitL_exit_CALC_SOFTMAX_LOOP_sva,
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_nl, COMPUTE_OUTER_LOOP_and_16_nl);
  assign CALC_EXP_LOOP_i_CALC_EXP_LOOP_i_nor_nl = ~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_1
      | (fsm_output[3]));
  assign CALC_EXP_LOOP_i_and_1_nl = lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_st_1_1
      & (~ (fsm_output[3]));
  assign CALC_SOFTMAX_LOOP_mux1h_22_nl = MUX1HOT_s_1_3_2(CALC_SOFTMAX_LOOP_equal_tmp_44_mx1w0,
      CALC_SOFTMAX_LOOP_equal_tmp_40_mx1w1, CALC_EXP_LOOP_and_svs_mx1w2, {and_dcpl_114
      , and_dcpl_115 , or_dcpl_6});
  assign COMPUTE_OUTER_LOOP_s_and_nl = (~ (fsm_output[1])) & or_tmp_47;
  assign COMPUTE_OUTER_LOOP_s_and_2_nl = (~ or_173_tmp) & (fsm_output[2]);
  assign COMPUTE_OUTER_LOOP_s_or_nl = (or_173_tmp & (fsm_output[2])) | (fsm_output[3]);
  assign or_269_nl = (fsm_output[4:2]!=3'b000);
  assign CALC_SOFTMAX_LOOP_mux_14_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_32_2,
      CALC_SOFTMAX_LOOP_equal_tmp_64_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_16_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_31_2,
      CALC_SOFTMAX_LOOP_equal_tmp_63_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_18_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_30_2,
      CALC_SOFTMAX_LOOP_equal_tmp_62_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_20_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_29_2,
      CALC_SOFTMAX_LOOP_equal_tmp_6_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_22_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_28_2,
      CALC_SOFTMAX_LOOP_equal_tmp_5_1, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_24_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_27_2,
      CALC_SOFTMAX_LOOP_equal_tmp_4_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_26_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_26_2,
      CALC_SOFTMAX_LOOP_equal_tmp_32_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_28_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_25_2,
      CALC_SOFTMAX_LOOP_equal_tmp_31_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_30_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_24_2,
      CALC_SOFTMAX_LOOP_equal_tmp_30_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_32_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_23_2,
      CALC_SOFTMAX_LOOP_equal_tmp_3_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_34_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_22_2,
      CALC_SOFTMAX_LOOP_equal_tmp_29_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_36_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_21_2,
      CALC_SOFTMAX_LOOP_equal_tmp_28_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_38_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_20_2,
      CALC_SOFTMAX_LOOP_equal_tmp_27_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_40_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_19_2,
      CALC_SOFTMAX_LOOP_equal_tmp_26_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_42_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_18_2,
      CALC_SOFTMAX_LOOP_equal_tmp_25_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_44_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_17_2,
      CALC_SOFTMAX_LOOP_equal_tmp_24_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_46_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_16_2,
      CALC_SOFTMAX_LOOP_equal_tmp_23_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_48_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_15_2,
      CALC_SOFTMAX_LOOP_equal_tmp_22_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_50_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_14_2,
      CALC_SOFTMAX_LOOP_equal_tmp_21_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_52_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_13_2,
      CALC_SOFTMAX_LOOP_equal_tmp_20_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_54_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_12_2,
      CALC_SOFTMAX_LOOP_equal_tmp_2_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_56_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_11_2,
      CALC_SOFTMAX_LOOP_equal_tmp_19_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_58_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_10_2,
      CALC_SOFTMAX_LOOP_equal_tmp_18_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_60_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_3_2,
      CALC_SOFTMAX_LOOP_equal_tmp_11_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_62_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_2_2,
      CALC_SOFTMAX_LOOP_equal_tmp_10_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_64_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_64_2,
      CALC_SOFTMAX_LOOP_equal_tmp_17_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_66_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_63_2,
      CALC_SOFTMAX_LOOP_equal_tmp_16_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_68_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_62_2,
      CALC_SOFTMAX_LOOP_equal_tmp_15_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_70_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_6_2,
      CALC_SOFTMAX_LOOP_equal_tmp_14_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_72_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_5_1,
      CALC_SOFTMAX_LOOP_equal_tmp_13_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign CALC_SOFTMAX_LOOP_mux_74_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_4_2,
      CALC_SOFTMAX_LOOP_equal_tmp_12_2, CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm_2);
  assign COMPUTE_OUTER_LOOP_mux_32_nl = MUX_s_1_2_2(exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_1,
      COMPUTE_OUTER_LOOP_stage_0_5, fsm_output[3]);
  assign COMPUTE_BATCH_LOOP_b_mux_nl = MUX_v_32_2_2(COMPUTE_BATCH_LOOP_b_sva, z_out_1,
      fsm_output[4]);
  assign softmax_softmax_not_nl = ~ (fsm_output[1]);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_4_nl = ~(CALC_SOFTMAX_LOOP_equal_tmp_66
      | CALC_SOFTMAX_LOOP_equal_tmp_67 | exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_1);
  assign CALC_SOFTMAX_LOOP_and_10_nl = CALC_EXP_LOOP_and_svs_mx1w2 & (~(CALC_SOFTMAX_LOOP_equal_tmp_66
      | CALC_SOFTMAX_LOOP_equal_tmp_67)) & (~ exit_COMPUTE_OUTER_LOOP_lpi_2_dfm_1);
  assign CALC_SOFTMAX_LOOP_mux_164_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_46_mx1w0,
      CALC_SOFTMAX_LOOP_equal_tmp_44_mx1w0, mux_tmp_35);
  assign CALC_SOFTMAX_LOOP_mux_166_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_47_mx1w0,
      CALC_SOFTMAX_LOOP_equal_tmp_46_mx1w0, mux_tmp_35);
  assign CALC_SOFTMAX_LOOP_mux_168_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_48_mx1w0,
      CALC_SOFTMAX_LOOP_equal_tmp_47_mx1w0, mux_tmp_35);
  assign CALC_SOFTMAX_LOOP_mux_170_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_equal_tmp_52_mx1w0,
      CALC_SOFTMAX_LOOP_equal_tmp_48_mx1w0, mux_tmp_35);
  assign CALC_SOFTMAX_LOOP_mux1h_228_nl = MUX1HOT_s_1_3_2(CALC_SOFTMAX_LOOP_nor_26_itm_mx1w0,
      CALC_SOFTMAX_LOOP_nor_32_itm_mx1w1, (CALC_EXP_LOOP_i_7_0_lpi_2_dfm_1_6_0_mx1[5]),
      {and_dcpl_114 , and_dcpl_115 , or_dcpl_6});
  assign nl_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_qif_acc_itm  =
      ({1'b1 , (~ libraries_leading_sign_74_0_5d32be77710879fd6707bb2fa0416553bf16_1)})
      + 8'b00110111;
  assign nor_nl = ~((CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[5]) | CALC_SOFTMAX_LOOP_slc_CALC_SOFTMAX_LOOP_i_7_0_6_5_itm);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_41_nl = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[3])
      & CALC_SOFTMAX_LOOP_nor_1_itm;
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_4_nl = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[1])
      & CALC_SOFTMAX_LOOP_nor_1_itm;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_nl
      = ~((SUM_EXP_LOOP_acc_1_tmp!=74'b00000000000000000000000000000000000000000000000000000000000000000000000000));
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_10_nl = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[3])
      & CALC_SOFTMAX_LOOP_nor_26_itm;
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_and_35_nl = (CALC_SOFTMAX_LOOP_i_7_0_lpi_2_6_0[1])
      & CALC_SOFTMAX_LOOP_nor_26_itm;
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_mux_68_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_asn_itm_1,
      CALC_SOFTMAX_LOOP_equal_tmp_42_mx1w2, lfst_exit_CALC_SOFTMAX_LOOP_lpi_2_dfm_1_1);
  assign COMPUTE_BATCH_LOOP_mux_4_nl = MUX_v_32_2_2((~ (conf_info[63:32])), z_out_1,
      fsm_output[4]);
  assign COMPUTE_BATCH_LOOP_or_1_nl = (~ (fsm_output[1])) | (fsm_output[4]);
  assign COMPUTE_BATCH_LOOP_mux_5_nl = MUX_v_32_2_2(32'b00000000000000000000000000000001,
      (~ (conf_info_crt_1_sva[63:32])), fsm_output[4]);
  assign nl_acc_nl = ({1'b1 , COMPUTE_BATCH_LOOP_mux_4_nl , COMPUTE_BATCH_LOOP_or_1_nl})
      + conv_u2u_33_34({COMPUTE_BATCH_LOOP_mux_5_nl , 1'b1});
  assign acc_nl = nl_acc_nl[33:0];
  assign z_out_32 = readslicef_34_1_33(acc_nl);
  assign COMPUTE_OUTER_LOOP_mux_34_nl = MUX_v_32_2_2(({7'b0000000 , COMPUTE_OUTER_LOOP_s_31_7_sva}),
      COMPUTE_BATCH_LOOP_b_sva, fsm_output[4]);
  assign nl_z_out_1 = COMPUTE_OUTER_LOOP_mux_34_nl + conv_s2u_2_32({(~ (fsm_output[4]))
      , 1'b1});
  assign z_out_1 = nl_z_out_1[31:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [24:0] MUX1HOT_v_25_4_2;
    input [24:0] input_3;
    input [24:0] input_2;
    input [24:0] input_1;
    input [24:0] input_0;
    input [3:0] sel;
    reg [24:0] result;
  begin
    result = input_0 & {25{sel[0]}};
    result = result | ( input_1 & {25{sel[1]}});
    result = result | ( input_2 & {25{sel[2]}});
    result = result | ( input_3 & {25{sel[3]}});
    MUX1HOT_v_25_4_2 = result;
  end
  endfunction


  function automatic [73:0] MUX1HOT_v_74_3_2;
    input [73:0] input_2;
    input [73:0] input_1;
    input [73:0] input_0;
    input [2:0] sel;
    reg [73:0] result;
  begin
    result = input_0 & {74{sel[0]}};
    result = result | ( input_1 & {74{sel[1]}});
    result = result | ( input_2 & {74{sel[2]}});
    MUX1HOT_v_74_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_8_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [9:0] input_2;
    input [9:0] input_3;
    input [9:0] input_4;
    input [9:0] input_5;
    input [9:0] input_6;
    input [9:0] input_7;
    input [2:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_10_8_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_32_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [31:0] input_3;
    input [31:0] input_4;
    input [31:0] input_5;
    input [31:0] input_6;
    input [31:0] input_7;
    input [31:0] input_8;
    input [31:0] input_9;
    input [31:0] input_10;
    input [31:0] input_11;
    input [31:0] input_12;
    input [31:0] input_13;
    input [31:0] input_14;
    input [31:0] input_15;
    input [31:0] input_16;
    input [31:0] input_17;
    input [31:0] input_18;
    input [31:0] input_19;
    input [31:0] input_20;
    input [31:0] input_21;
    input [31:0] input_22;
    input [31:0] input_23;
    input [31:0] input_24;
    input [31:0] input_25;
    input [31:0] input_26;
    input [31:0] input_27;
    input [31:0] input_28;
    input [31:0] input_29;
    input [31:0] input_30;
    input [31:0] input_31;
    input [4:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      5'b11000 : begin
        result = input_24;
      end
      5'b11001 : begin
        result = input_25;
      end
      5'b11010 : begin
        result = input_26;
      end
      5'b11011 : begin
        result = input_27;
      end
      5'b11100 : begin
        result = input_28;
      end
      5'b11101 : begin
        result = input_29;
      end
      5'b11110 : begin
        result = input_30;
      end
      default : begin
        result = input_31;
      end
    endcase
    MUX_v_32_32_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_4_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [1:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_3_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_4_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [4:0] input_2;
    input [4:0] input_3;
    input [1:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_5_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [73:0] MUX_v_74_2_2;
    input [73:0] input_0;
    input [73:0] input_1;
    input [0:0] sel;
    reg [73:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_74_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_4_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [6:0] input_2;
    input [6:0] input_3;
    input [1:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_7_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_8_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2 = result;
  end
  endfunction


  function automatic [93:0] MUX_v_94_2_2;
    input [93:0] input_0;
    input [93:0] input_1;
    input [0:0] sel;
    reg [93:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_94_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_34_1_33;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 33;
    readslicef_34_1_33 = tmp[0:0];
  end
  endfunction


  function automatic [18:0] readslicef_47_19_28;
    input [46:0] vector;
    reg [46:0] tmp;
  begin
    tmp = vector >> 28;
    readslicef_47_19_28 = tmp[18:0];
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input [0:0] vector;
  begin
    signext_7_1= {{6{vector[0]}}, vector};
  end
  endfunction


  function automatic [31:0] conv_s2u_2_32 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_32 = {{30{vector[1]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_s2u_9_11 = {{2{vector[8]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_11 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [18:0] conv_u2u_19_19 ;
    input [18:0]  vector ;
  begin
    conv_u2u_19_19 = vector;
  end
  endfunction


  function automatic [33:0] conv_u2u_33_34 ;
    input [32:0]  vector ;
  begin
    conv_u2u_33_34 = {1'b0, vector};
  end
  endfunction


  function automatic [73:0] conv_u2u_67_74 ;
    input [66:0]  vector ;
  begin
    conv_u2u_67_74 = {{7{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input_load_input
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input_load_input (
  clk, rst, conf_info, dma_read_ctrl_val, dma_read_ctrl_rdy, dma_read_ctrl_msg, dma_read_chnl_val,
      dma_read_chnl_rdy, dma_read_chnl_msg, done, input_ready_channel_val, input_ready_channel_rdy,
      input_ready_channel_msg, plm_in_cns_dat, plm_in_cns_vld, plm_in_cns_rdy, LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_clken_d,
      LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_d_d, LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d,
      LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_radr_d, LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_wadr_d,
      LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_we_d_pff
);
  input clk;
  input rst;
  input [63:0] conf_info;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  input done;
  input input_ready_channel_val;
  output input_ready_channel_rdy;
  input input_ready_channel_msg;
  output [4095:0] plm_in_cns_dat;
  output plm_in_cns_vld;
  input plm_in_cns_rdy;
  output LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_clken_d;
  output [31:0] LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_d_d;
  input [31:0] LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
  output [6:0] LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_radr_d;
  output [6:0] LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_wadr_d;
  output LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_we_d_pff;


  // Interconnect Declarations
  wire load_input_wen;
  wire dma_read_ctrl_Push_mioi_wen_comp;
  wire dma_read_chnl_Pop_mioi_wen_comp;
  wire [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt;
  wire input_ready_channel_Pop_mioi_wen_comp;
  wire plm_in_cnsi_wen_comp;
  reg [31:0] plm_in_cnsi_idat_4095_4064;
  reg [31:0] plm_in_cnsi_idat_4063_4032;
  reg [31:0] plm_in_cnsi_idat_4031_4000;
  reg [31:0] plm_in_cnsi_idat_3999_3968;
  reg [31:0] plm_in_cnsi_idat_3967_3936;
  reg [31:0] plm_in_cnsi_idat_3935_3904;
  reg [31:0] plm_in_cnsi_idat_3903_3872;
  reg [31:0] plm_in_cnsi_idat_3871_3840;
  reg [31:0] plm_in_cnsi_idat_3839_3808;
  reg [31:0] plm_in_cnsi_idat_3807_3776;
  reg [31:0] plm_in_cnsi_idat_3775_3744;
  reg [31:0] plm_in_cnsi_idat_3743_3712;
  reg [31:0] plm_in_cnsi_idat_3711_3680;
  reg [31:0] plm_in_cnsi_idat_3679_3648;
  reg [31:0] plm_in_cnsi_idat_3647_3616;
  reg [31:0] plm_in_cnsi_idat_3615_3584;
  reg [31:0] plm_in_cnsi_idat_3583_3552;
  reg [31:0] plm_in_cnsi_idat_3551_3520;
  reg [31:0] plm_in_cnsi_idat_3519_3488;
  reg [31:0] plm_in_cnsi_idat_3487_3456;
  reg [31:0] plm_in_cnsi_idat_3455_3424;
  reg [31:0] plm_in_cnsi_idat_3423_3392;
  reg [31:0] plm_in_cnsi_idat_3391_3360;
  reg [31:0] plm_in_cnsi_idat_3359_3328;
  reg [31:0] plm_in_cnsi_idat_3327_3296;
  reg [31:0] plm_in_cnsi_idat_3295_3264;
  reg [31:0] plm_in_cnsi_idat_3263_3232;
  reg [31:0] plm_in_cnsi_idat_3231_3200;
  reg [31:0] plm_in_cnsi_idat_3199_3168;
  reg [31:0] plm_in_cnsi_idat_3167_3136;
  reg [31:0] plm_in_cnsi_idat_3135_3104;
  reg [31:0] plm_in_cnsi_idat_3103_3072;
  reg [31:0] plm_in_cnsi_idat_3071_3040;
  reg [31:0] plm_in_cnsi_idat_3039_3008;
  reg [31:0] plm_in_cnsi_idat_3007_2976;
  reg [31:0] plm_in_cnsi_idat_2975_2944;
  reg [31:0] plm_in_cnsi_idat_2943_2912;
  reg [31:0] plm_in_cnsi_idat_2911_2880;
  reg [31:0] plm_in_cnsi_idat_2879_2848;
  reg [31:0] plm_in_cnsi_idat_2847_2816;
  reg [31:0] plm_in_cnsi_idat_2815_2784;
  reg [31:0] plm_in_cnsi_idat_2783_2752;
  reg [31:0] plm_in_cnsi_idat_2751_2720;
  reg [31:0] plm_in_cnsi_idat_2719_2688;
  reg [31:0] plm_in_cnsi_idat_2687_2656;
  reg [31:0] plm_in_cnsi_idat_2655_2624;
  reg [31:0] plm_in_cnsi_idat_2623_2592;
  reg [31:0] plm_in_cnsi_idat_2591_2560;
  reg [31:0] plm_in_cnsi_idat_2559_2528;
  reg [31:0] plm_in_cnsi_idat_2527_2496;
  reg [31:0] plm_in_cnsi_idat_2495_2464;
  reg [31:0] plm_in_cnsi_idat_2463_2432;
  reg [31:0] plm_in_cnsi_idat_2431_2400;
  reg [31:0] plm_in_cnsi_idat_2399_2368;
  reg [31:0] plm_in_cnsi_idat_2367_2336;
  reg [31:0] plm_in_cnsi_idat_2335_2304;
  reg [31:0] plm_in_cnsi_idat_2303_2272;
  reg [31:0] plm_in_cnsi_idat_2271_2240;
  reg [31:0] plm_in_cnsi_idat_2239_2208;
  reg [31:0] plm_in_cnsi_idat_2207_2176;
  reg [31:0] plm_in_cnsi_idat_2175_2144;
  reg [31:0] plm_in_cnsi_idat_2143_2112;
  reg [31:0] plm_in_cnsi_idat_2111_2080;
  reg [31:0] plm_in_cnsi_idat_2079_2048;
  reg [31:0] plm_in_cnsi_idat_2047_2016;
  reg [31:0] plm_in_cnsi_idat_2015_1984;
  reg [31:0] plm_in_cnsi_idat_1983_1952;
  reg [31:0] plm_in_cnsi_idat_1951_1920;
  reg [31:0] plm_in_cnsi_idat_1919_1888;
  reg [31:0] plm_in_cnsi_idat_1887_1856;
  reg [31:0] plm_in_cnsi_idat_1855_1824;
  reg [31:0] plm_in_cnsi_idat_1823_1792;
  reg [31:0] plm_in_cnsi_idat_1791_1760;
  reg [31:0] plm_in_cnsi_idat_1759_1728;
  reg [31:0] plm_in_cnsi_idat_1727_1696;
  reg [31:0] plm_in_cnsi_idat_1695_1664;
  reg [31:0] plm_in_cnsi_idat_1663_1632;
  reg [31:0] plm_in_cnsi_idat_1631_1600;
  reg [31:0] plm_in_cnsi_idat_1599_1568;
  reg [31:0] plm_in_cnsi_idat_1567_1536;
  reg [31:0] plm_in_cnsi_idat_1535_1504;
  reg [31:0] plm_in_cnsi_idat_1503_1472;
  reg [31:0] plm_in_cnsi_idat_1471_1440;
  reg [31:0] plm_in_cnsi_idat_1439_1408;
  reg [31:0] plm_in_cnsi_idat_1407_1376;
  reg [31:0] plm_in_cnsi_idat_1375_1344;
  reg [31:0] plm_in_cnsi_idat_1343_1312;
  reg [31:0] plm_in_cnsi_idat_1311_1280;
  reg [31:0] plm_in_cnsi_idat_1279_1248;
  reg [31:0] plm_in_cnsi_idat_1247_1216;
  reg [31:0] plm_in_cnsi_idat_1215_1184;
  reg [31:0] plm_in_cnsi_idat_1183_1152;
  reg [31:0] plm_in_cnsi_idat_1151_1120;
  reg [31:0] plm_in_cnsi_idat_1119_1088;
  reg [31:0] plm_in_cnsi_idat_1087_1056;
  reg [31:0] plm_in_cnsi_idat_1055_1024;
  reg [31:0] plm_in_cnsi_idat_1023_992;
  reg [31:0] plm_in_cnsi_idat_991_960;
  reg [31:0] plm_in_cnsi_idat_959_928;
  reg [31:0] plm_in_cnsi_idat_927_896;
  reg [31:0] plm_in_cnsi_idat_895_864;
  reg [31:0] plm_in_cnsi_idat_863_832;
  reg [31:0] plm_in_cnsi_idat_831_800;
  reg [31:0] plm_in_cnsi_idat_799_768;
  reg [31:0] plm_in_cnsi_idat_767_736;
  reg [31:0] plm_in_cnsi_idat_735_704;
  reg [31:0] plm_in_cnsi_idat_703_672;
  reg [31:0] plm_in_cnsi_idat_671_640;
  reg [31:0] plm_in_cnsi_idat_639_608;
  reg [31:0] plm_in_cnsi_idat_607_576;
  reg [31:0] plm_in_cnsi_idat_575_544;
  reg [31:0] plm_in_cnsi_idat_543_512;
  reg [31:0] plm_in_cnsi_idat_511_480;
  reg [31:0] plm_in_cnsi_idat_479_448;
  reg [31:0] plm_in_cnsi_idat_447_416;
  reg [31:0] plm_in_cnsi_idat_415_384;
  reg [31:0] plm_in_cnsi_idat_383_352;
  reg [31:0] plm_in_cnsi_idat_351_320;
  reg [31:0] plm_in_cnsi_idat_319_288;
  reg [31:0] plm_in_cnsi_idat_287_256;
  reg [31:0] plm_in_cnsi_idat_255_224;
  reg [31:0] plm_in_cnsi_idat_223_192;
  reg [31:0] plm_in_cnsi_idat_191_160;
  reg [31:0] plm_in_cnsi_idat_159_128;
  reg [31:0] plm_in_cnsi_idat_127_96;
  reg [31:0] plm_in_cnsi_idat_95_64;
  reg [31:0] plm_in_cnsi_idat_63_32;
  reg [31:0] plm_in_cnsi_idat_31_0;
  wire [7:0] fsm_output;
  wire or_tmp_4;
  wire and_tmp;
  wire mux_tmp_2;
  wire mux_tmp_3;
  wire mux_tmp_4;
  wire mux_tmp_5;
  wire mux_tmp_8;
  wire and_dcpl_7;
  wire and_dcpl_8;
  wire and_dcpl_9;
  wire and_dcpl_10;
  wire and_dcpl_11;
  wire and_dcpl_13;
  wire and_dcpl_14;
  wire and_dcpl_15;
  wire and_dcpl_17;
  wire and_dcpl_18;
  wire and_dcpl_20;
  wire and_dcpl_21;
  wire and_dcpl_23;
  wire and_dcpl_25;
  wire and_dcpl_26;
  wire and_dcpl_28;
  wire and_dcpl_30;
  wire and_dcpl_32;
  wire and_dcpl_34;
  wire and_dcpl_35;
  wire and_dcpl_36;
  wire and_dcpl_37;
  wire and_dcpl_39;
  wire and_dcpl_41;
  wire and_dcpl_43;
  wire and_dcpl_45;
  wire and_dcpl_47;
  wire and_dcpl_49;
  wire and_dcpl_60;
  wire and_dcpl_61;
  wire and_dcpl_78;
  wire and_dcpl_95;
  wire and_dcpl_96;
  wire and_dcpl_113;
  wire and_dcpl_130;
  wire and_dcpl_131;
  wire and_dcpl_148;
  wire and_dcpl_166;
  wire and_dcpl_170;
  wire and_dcpl_175;
  wire and_dcpl_179;
  wire or_dcpl_5;
  wire or_dcpl_6;
  wire or_dcpl_7;
  wire or_dcpl_9;
  wire and_dcpl_187;
  wire and_dcpl_188;
  wire and_dcpl_189;
  wire or_dcpl_21;
  wire or_dcpl_22;
  wire or_dcpl_23;
  wire or_dcpl_24;
  wire or_dcpl_25;
  wire and_dcpl_202;
  wire or_dcpl_32;
  wire or_dcpl_34;
  wire or_dcpl_35;
  wire or_dcpl_36;
  wire or_dcpl_38;
  wire or_dcpl_39;
  wire or_dcpl_41;
  wire or_dcpl_43;
  wire or_dcpl_45;
  wire or_dcpl_46;
  wire or_dcpl_48;
  wire or_dcpl_50;
  wire or_dcpl_52;
  wire or_dcpl_54;
  wire or_dcpl_55;
  wire or_dcpl_56;
  wire or_dcpl_58;
  wire or_dcpl_60;
  wire or_dcpl_63;
  wire or_dcpl_65;
  wire or_dcpl_77;
  wire or_dcpl_78;
  wire or_dcpl_95;
  wire or_dcpl_112;
  wire or_dcpl_113;
  wire or_dcpl_130;
  wire or_dcpl_147;
  wire or_dcpl_148;
  wire or_dcpl_165;
  reg LOAD_DATA_INNER_LOOP_stage_0;
  reg LOAD_DATA_INNER_LOOP_stage_0_2;
  reg exit_LOAD_DATA_INNER_LOOP_sva_st_1;
  wire and_205_cse;
  reg reg_dma_read_ctrl_Push_mioi_oswt_cse;
  reg reg_dma_read_chnl_Pop_mioi_oswt_cse;
  reg reg_input_ready_channel_Pop_mioi_oswt_cse;
  wire LOAD_DATA_OUTER_LOOP_and_cse;
  wire or_8_cse;
  wire or_11_cse;
  wire nor_6_cse;
  wire mux_4_cse;
  wire or_1_cse;
  wire and_183_rmff;
  wire and_186_rmff;
  wire and_187_rmff;
  reg [31:0] offset_lpi_2;
  reg [24:0] LOAD_DATA_OUTER_LOOP_s_31_7_sva;
  wire [6:0] LOAD_DATA_OUTER_LOOP_len_qr_6_0_lpi_2_dfm_1;
  reg [6:0] LOAD_DATA_INNER_LOOP_slc_LOAD_DATA_INNER_LOOP_i_6_0_itm_1;
  wire and_dcpl_214;
  wire [31:0] z_out;
  wire [32:0] nl_z_out;
  wire and_dcpl_215;
  wire and_dcpl_216;
  wire and_dcpl_219;
  wire and_dcpl_220;
  wire and_dcpl_221;
  wire and_dcpl_222;
  wire and_dcpl_227;
  wire and_dcpl_228;
  wire and_dcpl_230;
  wire and_dcpl_233;
  wire and_dcpl_235;
  wire and_dcpl_238;
  wire and_dcpl_249;
  wire [24:0] z_out_2;
  wire [25:0] nl_z_out_2;
  reg [63:0] conf_info_crt_sva;
  reg [31:0] LOAD_BATCH_LOOP_b_sva;
  reg [6:0] LOAD_DATA_OUTER_LOOP_len_qr_6_0_lpi_2_dfm;
  reg [15:0] LOAD_DATA_INNER_LOOP_i_sva;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_8_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_9_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_10_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_11_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_12_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_13_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_14_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_15_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_16_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_17_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_18_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_19_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_20_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_21_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_22_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_23_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_24_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_25_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_26_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_27_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_28_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_29_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_30_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_31_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_32_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_33_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_34_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_35_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_36_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_37_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_38_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_39_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_40_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_41_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_42_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_43_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_44_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_45_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_46_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_47_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_48_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_49_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_50_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_51_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_52_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_53_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_54_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_55_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_56_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_57_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_58_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_59_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_60_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_61_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_62_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_63_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_64_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_65_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_66_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_67_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_68_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_69_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_70_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_71_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_72_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_73_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_74_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_75_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_76_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_77_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_78_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_79_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_80_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_81_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_82_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_83_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_84_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_85_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_86_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_87_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_88_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_89_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_90_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_91_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_92_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_93_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_94_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_95_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_96_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_97_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_98_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_99_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_100_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_101_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_102_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_103_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_104_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_105_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_106_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_107_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_108_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_109_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_110_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_111_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_112_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_113_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_114_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_115_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_116_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_117_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_118_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_119_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_120_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_121_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_122_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_123_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_124_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_125_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_126_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_127_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_128_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_129_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_130_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_131_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_132_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_133_itm;
  reg [31:0] LOAD_DATA_OUTER_LOOP_asn_134_itm;
  wire LOAD_DATA_INNER_LOOP_stage_0_mx0c0;
  wire LOAD_BATCH_LOOP_or_1_ssc;
  wire nor_16_cse;
  wire z_out_1_32;

  wire[0:0] mux_35_nl;
  wire[0:0] mux_13_nl;
  wire[31:0] LOAD_BATCH_LOOP_b_mux_nl;
  wire[0:0] mux_21_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] mux_37_nl;
  wire[0:0] not_nl;
  wire[0:0] and_192_nl;
  wire[0:0] mux_42_nl;
  wire[0:0] mux_41_nl;
  wire[0:0] nor_3_nl;
  wire[24:0] LOAD_DATA_OUTER_LOOP_len_qif_mux1h_nl;
  wire[0:0] or_37_nl;
  wire[0:0] mux_44_nl;
  wire[0:0] nor_4_nl;
  wire[0:0] and_196_nl;
  wire[0:0] and_198_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] LOAD_DATA_OUTER_LOOP_mux_nl;
  wire[0:0] dma_read_ctrl_write_reset_check_ResetChecker_dma_read_ctrl_write_reset_check_ResetChecker_and_nl;
  wire[0:0] LOAD_DATA_OUTER_LOOP_len_not_4_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] mux_10_nl;
  wire[6:0] nor_12_nl;
  wire[6:0] mux1h_nl;
  wire[0:0] and_13_nl;
  wire[0:0] and_17_nl;
  wire[0:0] and_20_nl;
  wire[0:0] and_23_nl;
  wire[0:0] and_25_nl;
  wire[0:0] and_28_nl;
  wire[0:0] and_30_nl;
  wire[0:0] and_32_nl;
  wire[0:0] and_34_nl;
  wire[0:0] and_39_nl;
  wire[0:0] and_41_nl;
  wire[0:0] and_43_nl;
  wire[0:0] and_45_nl;
  wire[0:0] and_47_nl;
  wire[0:0] and_49_nl;
  wire[0:0] and_51_nl;
  wire[0:0] and_52_nl;
  wire[0:0] and_53_nl;
  wire[0:0] and_54_nl;
  wire[0:0] and_55_nl;
  wire[0:0] and_56_nl;
  wire[0:0] and_57_nl;
  wire[0:0] and_58_nl;
  wire[0:0] and_59_nl;
  wire[0:0] and_60_nl;
  wire[0:0] and_63_nl;
  wire[0:0] and_64_nl;
  wire[0:0] and_65_nl;
  wire[0:0] and_66_nl;
  wire[0:0] and_67_nl;
  wire[0:0] and_68_nl;
  wire[0:0] and_69_nl;
  wire[0:0] and_70_nl;
  wire[0:0] and_71_nl;
  wire[0:0] and_72_nl;
  wire[0:0] and_73_nl;
  wire[0:0] and_74_nl;
  wire[0:0] and_75_nl;
  wire[0:0] and_76_nl;
  wire[0:0] and_77_nl;
  wire[0:0] and_78_nl;
  wire[0:0] and_80_nl;
  wire[0:0] and_81_nl;
  wire[0:0] and_82_nl;
  wire[0:0] and_83_nl;
  wire[0:0] and_84_nl;
  wire[0:0] and_85_nl;
  wire[0:0] and_86_nl;
  wire[0:0] and_87_nl;
  wire[0:0] and_88_nl;
  wire[0:0] and_89_nl;
  wire[0:0] and_90_nl;
  wire[0:0] and_91_nl;
  wire[0:0] and_92_nl;
  wire[0:0] and_93_nl;
  wire[0:0] and_94_nl;
  wire[0:0] and_95_nl;
  wire[0:0] and_98_nl;
  wire[0:0] and_99_nl;
  wire[0:0] and_100_nl;
  wire[0:0] and_101_nl;
  wire[0:0] and_102_nl;
  wire[0:0] and_103_nl;
  wire[0:0] and_104_nl;
  wire[0:0] and_105_nl;
  wire[0:0] and_106_nl;
  wire[0:0] and_107_nl;
  wire[0:0] and_108_nl;
  wire[0:0] and_109_nl;
  wire[0:0] and_110_nl;
  wire[0:0] and_111_nl;
  wire[0:0] and_112_nl;
  wire[0:0] and_113_nl;
  wire[0:0] and_115_nl;
  wire[0:0] and_116_nl;
  wire[0:0] and_117_nl;
  wire[0:0] and_118_nl;
  wire[0:0] and_119_nl;
  wire[0:0] and_120_nl;
  wire[0:0] and_121_nl;
  wire[0:0] and_122_nl;
  wire[0:0] and_123_nl;
  wire[0:0] and_124_nl;
  wire[0:0] and_125_nl;
  wire[0:0] and_126_nl;
  wire[0:0] and_127_nl;
  wire[0:0] and_128_nl;
  wire[0:0] and_129_nl;
  wire[0:0] and_130_nl;
  wire[0:0] and_133_nl;
  wire[0:0] and_134_nl;
  wire[0:0] and_135_nl;
  wire[0:0] and_136_nl;
  wire[0:0] and_137_nl;
  wire[0:0] and_138_nl;
  wire[0:0] and_139_nl;
  wire[0:0] and_140_nl;
  wire[0:0] and_141_nl;
  wire[0:0] and_142_nl;
  wire[0:0] and_143_nl;
  wire[0:0] and_144_nl;
  wire[0:0] and_145_nl;
  wire[0:0] and_146_nl;
  wire[0:0] and_147_nl;
  wire[0:0] and_148_nl;
  wire[0:0] and_150_nl;
  wire[0:0] and_151_nl;
  wire[0:0] and_152_nl;
  wire[0:0] and_153_nl;
  wire[0:0] and_154_nl;
  wire[0:0] and_155_nl;
  wire[0:0] and_156_nl;
  wire[0:0] and_157_nl;
  wire[0:0] and_158_nl;
  wire[0:0] and_159_nl;
  wire[0:0] and_160_nl;
  wire[0:0] and_161_nl;
  wire[0:0] and_162_nl;
  wire[0:0] and_163_nl;
  wire[0:0] and_164_nl;
  wire[0:0] and_165_nl;
  wire[0:0] and_168_nl;
  wire[0:0] and_169_nl;
  wire[0:0] and_170_nl;
  wire[0:0] and_172_nl;
  wire[0:0] mux_28_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] mux_25_nl;
  wire[0:0] or_12_nl;
  wire[0:0] mux_24_nl;
  wire[0:0] or_9_nl;
  wire[0:0] and_173_nl;
  wire[31:0] LOAD_DATA_OUTER_LOOP_mux_131_nl;
  wire[24:0] LOAD_DATA_OUTER_LOOP_LOAD_DATA_OUTER_LOOP_and_1_nl;
  wire[0:0] not_116_nl;
  wire[6:0] LOAD_DATA_OUTER_LOOP_mux_132_nl;
  wire[33:0] acc_1_nl;
  wire[34:0] nl_acc_1_nl;
  wire[31:0] LOAD_BATCH_LOOP_mux1h_3_nl;
  wire[0:0] LOAD_BATCH_LOOP_or_2_nl;
  wire[24:0] LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_nor_1_nl;
  wire[24:0] LOAD_BATCH_LOOP_mux1h_4_nl;
  wire[6:0] LOAD_BATCH_LOOP_mux1h_5_nl;
  wire[24:0] LOAD_DATA_INNER_LOOP_mux_127_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input;
  assign nl_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input
      = offset_lpi_2;
  wire[24:0] LOAD_DATA_OUTER_LOOP_len_qif_mux_nl;
  wire [31:0] nl_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_length_rsc_dat_load_input;
  assign LOAD_DATA_OUTER_LOOP_len_qif_mux_nl = MUX_v_25_2_2(LOAD_DATA_OUTER_LOOP_s_31_7_sva,
      25'b0000000000000000000000001, z_out_1_32);
  assign nl_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_length_rsc_dat_load_input
      = {LOAD_DATA_OUTER_LOOP_len_qif_mux_nl , LOAD_DATA_OUTER_LOOP_len_qr_6_0_lpi_2_dfm_1};
  wire [4095:0] nl_softmax_load_input_load_input_plm_in_cnsi_inst_plm_in_cnsi_idat;
  assign nl_softmax_load_input_load_input_plm_in_cnsi_inst_plm_in_cnsi_idat = {plm_in_cnsi_idat_4095_4064
      , plm_in_cnsi_idat_4063_4032 , plm_in_cnsi_idat_4031_4000 , plm_in_cnsi_idat_3999_3968
      , plm_in_cnsi_idat_3967_3936 , plm_in_cnsi_idat_3935_3904 , plm_in_cnsi_idat_3903_3872
      , plm_in_cnsi_idat_3871_3840 , plm_in_cnsi_idat_3839_3808 , plm_in_cnsi_idat_3807_3776
      , plm_in_cnsi_idat_3775_3744 , plm_in_cnsi_idat_3743_3712 , plm_in_cnsi_idat_3711_3680
      , plm_in_cnsi_idat_3679_3648 , plm_in_cnsi_idat_3647_3616 , plm_in_cnsi_idat_3615_3584
      , plm_in_cnsi_idat_3583_3552 , plm_in_cnsi_idat_3551_3520 , plm_in_cnsi_idat_3519_3488
      , plm_in_cnsi_idat_3487_3456 , plm_in_cnsi_idat_3455_3424 , plm_in_cnsi_idat_3423_3392
      , plm_in_cnsi_idat_3391_3360 , plm_in_cnsi_idat_3359_3328 , plm_in_cnsi_idat_3327_3296
      , plm_in_cnsi_idat_3295_3264 , plm_in_cnsi_idat_3263_3232 , plm_in_cnsi_idat_3231_3200
      , plm_in_cnsi_idat_3199_3168 , plm_in_cnsi_idat_3167_3136 , plm_in_cnsi_idat_3135_3104
      , plm_in_cnsi_idat_3103_3072 , plm_in_cnsi_idat_3071_3040 , plm_in_cnsi_idat_3039_3008
      , plm_in_cnsi_idat_3007_2976 , plm_in_cnsi_idat_2975_2944 , plm_in_cnsi_idat_2943_2912
      , plm_in_cnsi_idat_2911_2880 , plm_in_cnsi_idat_2879_2848 , plm_in_cnsi_idat_2847_2816
      , plm_in_cnsi_idat_2815_2784 , plm_in_cnsi_idat_2783_2752 , plm_in_cnsi_idat_2751_2720
      , plm_in_cnsi_idat_2719_2688 , plm_in_cnsi_idat_2687_2656 , plm_in_cnsi_idat_2655_2624
      , plm_in_cnsi_idat_2623_2592 , plm_in_cnsi_idat_2591_2560 , plm_in_cnsi_idat_2559_2528
      , plm_in_cnsi_idat_2527_2496 , plm_in_cnsi_idat_2495_2464 , plm_in_cnsi_idat_2463_2432
      , plm_in_cnsi_idat_2431_2400 , plm_in_cnsi_idat_2399_2368 , plm_in_cnsi_idat_2367_2336
      , plm_in_cnsi_idat_2335_2304 , plm_in_cnsi_idat_2303_2272 , plm_in_cnsi_idat_2271_2240
      , plm_in_cnsi_idat_2239_2208 , plm_in_cnsi_idat_2207_2176 , plm_in_cnsi_idat_2175_2144
      , plm_in_cnsi_idat_2143_2112 , plm_in_cnsi_idat_2111_2080 , plm_in_cnsi_idat_2079_2048
      , plm_in_cnsi_idat_2047_2016 , plm_in_cnsi_idat_2015_1984 , plm_in_cnsi_idat_1983_1952
      , plm_in_cnsi_idat_1951_1920 , plm_in_cnsi_idat_1919_1888 , plm_in_cnsi_idat_1887_1856
      , plm_in_cnsi_idat_1855_1824 , plm_in_cnsi_idat_1823_1792 , plm_in_cnsi_idat_1791_1760
      , plm_in_cnsi_idat_1759_1728 , plm_in_cnsi_idat_1727_1696 , plm_in_cnsi_idat_1695_1664
      , plm_in_cnsi_idat_1663_1632 , plm_in_cnsi_idat_1631_1600 , plm_in_cnsi_idat_1599_1568
      , plm_in_cnsi_idat_1567_1536 , plm_in_cnsi_idat_1535_1504 , plm_in_cnsi_idat_1503_1472
      , plm_in_cnsi_idat_1471_1440 , plm_in_cnsi_idat_1439_1408 , plm_in_cnsi_idat_1407_1376
      , plm_in_cnsi_idat_1375_1344 , plm_in_cnsi_idat_1343_1312 , plm_in_cnsi_idat_1311_1280
      , plm_in_cnsi_idat_1279_1248 , plm_in_cnsi_idat_1247_1216 , plm_in_cnsi_idat_1215_1184
      , plm_in_cnsi_idat_1183_1152 , plm_in_cnsi_idat_1151_1120 , plm_in_cnsi_idat_1119_1088
      , plm_in_cnsi_idat_1087_1056 , plm_in_cnsi_idat_1055_1024 , plm_in_cnsi_idat_1023_992
      , plm_in_cnsi_idat_991_960 , plm_in_cnsi_idat_959_928 , plm_in_cnsi_idat_927_896
      , plm_in_cnsi_idat_895_864 , plm_in_cnsi_idat_863_832 , plm_in_cnsi_idat_831_800
      , plm_in_cnsi_idat_799_768 , plm_in_cnsi_idat_767_736 , plm_in_cnsi_idat_735_704
      , plm_in_cnsi_idat_703_672 , plm_in_cnsi_idat_671_640 , plm_in_cnsi_idat_639_608
      , plm_in_cnsi_idat_607_576 , plm_in_cnsi_idat_575_544 , plm_in_cnsi_idat_543_512
      , plm_in_cnsi_idat_511_480 , plm_in_cnsi_idat_479_448 , plm_in_cnsi_idat_447_416
      , plm_in_cnsi_idat_415_384 , plm_in_cnsi_idat_383_352 , plm_in_cnsi_idat_351_320
      , plm_in_cnsi_idat_319_288 , plm_in_cnsi_idat_287_256 , plm_in_cnsi_idat_255_224
      , plm_in_cnsi_idat_223_192 , plm_in_cnsi_idat_191_160 , plm_in_cnsi_idat_159_128
      , plm_in_cnsi_idat_127_96 , plm_in_cnsi_idat_95_64 , plm_in_cnsi_idat_63_32
      , plm_in_cnsi_idat_31_0};
  wire [0:0] nl_softmax_load_input_load_input_load_input_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0;
  assign nl_softmax_load_input_load_input_load_input_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0
      = ~ done;
  wire [0:0] nl_softmax_load_input_load_input_load_input_fsm_inst_LOAD_BATCH_LOOP_C_0_tr0;
  assign nl_softmax_load_input_load_input_load_input_fsm_inst_LOAD_BATCH_LOOP_C_0_tr0
      = ~ z_out_1_32;
  wire [0:0] nl_softmax_load_input_load_input_load_input_fsm_inst_LOAD_DATA_INNER_LOOP_C_0_tr0;
  assign nl_softmax_load_input_load_input_load_input_fsm_inst_LOAD_DATA_INNER_LOOP_C_0_tr0
      = ~(LOAD_DATA_INNER_LOOP_stage_0 | LOAD_DATA_INNER_LOOP_stage_0_2);
  esp_acc_softmax_softmax_load_input_load_input_dma_read_ctrl_Push_mioi softmax_load_input_load_input_dma_read_ctrl_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_ctrl_val(dma_read_ctrl_val),
      .dma_read_ctrl_rdy(dma_read_ctrl_rdy),
      .dma_read_ctrl_msg(dma_read_ctrl_msg),
      .load_input_wen(load_input_wen),
      .dma_read_ctrl_Push_mioi_oswt(reg_dma_read_ctrl_Push_mioi_oswt_cse),
      .dma_read_ctrl_Push_mioi_wen_comp(dma_read_ctrl_Push_mioi_wen_comp),
      .dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input(nl_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat_load_input[31:0]),
      .dma_read_ctrl_Push_mioi_m_length_rsc_dat_load_input(nl_softmax_load_input_load_input_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_length_rsc_dat_load_input[31:0]),
      .dma_read_ctrl_Push_mioi_oswt_pff(and_183_rmff)
    );
  esp_acc_softmax_softmax_load_input_load_input_dma_read_chnl_Pop_mioi softmax_load_input_load_input_dma_read_chnl_Pop_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_chnl_val(dma_read_chnl_val),
      .dma_read_chnl_rdy(dma_read_chnl_rdy),
      .dma_read_chnl_msg(dma_read_chnl_msg),
      .load_input_wen(load_input_wen),
      .dma_read_chnl_Pop_mioi_oswt(reg_dma_read_chnl_Pop_mioi_oswt_cse),
      .dma_read_chnl_Pop_mioi_wen_comp(dma_read_chnl_Pop_mioi_wen_comp),
      .dma_read_chnl_Pop_mioi_return_rsc_z_mxwt(dma_read_chnl_Pop_mioi_return_rsc_z_mxwt),
      .dma_read_chnl_Pop_mioi_oswt_pff(and_186_rmff)
    );
  esp_acc_softmax_softmax_load_input_load_input_input_ready_channel_Pop_mioi softmax_load_input_load_input_input_ready_channel_Pop_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .input_ready_channel_val(input_ready_channel_val),
      .input_ready_channel_rdy(input_ready_channel_rdy),
      .input_ready_channel_msg(input_ready_channel_msg),
      .load_input_wen(load_input_wen),
      .input_ready_channel_Pop_mioi_oswt(reg_input_ready_channel_Pop_mioi_oswt_cse),
      .input_ready_channel_Pop_mioi_wen_comp(input_ready_channel_Pop_mioi_wen_comp),
      .input_ready_channel_Pop_mioi_oswt_pff(and_187_rmff)
    );
  esp_acc_softmax_softmax_load_input_load_input_plm_in_cnsi softmax_load_input_load_input_plm_in_cnsi_inst
      (
      .clk(clk),
      .rst(rst),
      .plm_in_cns_dat(plm_in_cns_dat),
      .plm_in_cns_vld(plm_in_cns_vld),
      .plm_in_cns_rdy(plm_in_cns_rdy),
      .load_input_wen(load_input_wen),
      .plm_in_cnsi_oswt(reg_input_ready_channel_Pop_mioi_oswt_cse),
      .plm_in_cnsi_wen_comp(plm_in_cnsi_wen_comp),
      .plm_in_cnsi_idat(nl_softmax_load_input_load_input_plm_in_cnsi_inst_plm_in_cnsi_idat[4095:0])
    );
  esp_acc_softmax_softmax_load_input_load_input_staller softmax_load_input_load_input_staller_inst
      (
      .load_input_wen(load_input_wen),
      .dma_read_ctrl_Push_mioi_wen_comp(dma_read_ctrl_Push_mioi_wen_comp),
      .dma_read_chnl_Pop_mioi_wen_comp(dma_read_chnl_Pop_mioi_wen_comp),
      .input_ready_channel_Pop_mioi_wen_comp(input_ready_channel_Pop_mioi_wen_comp),
      .plm_in_cnsi_wen_comp(plm_in_cnsi_wen_comp)
    );
  esp_acc_softmax_softmax_load_input_load_input_load_input_fsm softmax_load_input_load_input_load_input_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .load_input_wen(load_input_wen),
      .fsm_output(fsm_output),
      .WAIT_FOR_CONFIG_LOOP_C_0_tr0(nl_softmax_load_input_load_input_load_input_fsm_inst_WAIT_FOR_CONFIG_LOOP_C_0_tr0[0:0]),
      .load_input_rlp_C_0_tr0(z_out_1_32),
      .LOAD_BATCH_LOOP_C_0_tr0(nl_softmax_load_input_load_input_load_input_fsm_inst_LOAD_BATCH_LOOP_C_0_tr0[0:0]),
      .LOAD_DATA_INNER_LOOP_C_0_tr0(nl_softmax_load_input_load_input_load_input_fsm_inst_LOAD_DATA_INNER_LOOP_C_0_tr0[0:0]),
      .LOAD_DATA_OUTER_LOOP_C_131_tr0(LOAD_DATA_INNER_LOOP_stage_0),
      .LOAD_BATCH_LOOP_C_1_tr0(z_out_1_32)
    );
  assign LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_clken_d = load_input_wen;
  assign and_205_cse = (fsm_output[2:1]==2'b11);
  assign or_11_cse = (fsm_output[4:3]!=2'b00);
  assign and_183_rmff = and_dcpl_11 & and_dcpl_43;
  assign and_186_rmff = and_dcpl_179 & and_dcpl_175 & LOAD_DATA_INNER_LOOP_stage_0
      & z_out_1_32;
  assign and_187_rmff = and_dcpl_166 & and_dcpl_49;
  assign LOAD_DATA_OUTER_LOOP_and_cse = load_input_wen & (~(or_dcpl_9 | or_dcpl_7));
  assign or_8_cse = (fsm_output[2:1]!=2'b00);
  assign nor_6_cse = ~((fsm_output[4:3]!=2'b00));
  assign mux_4_cse = MUX_s_1_2_2((~ (fsm_output[2])), (fsm_output[2]), fsm_output[1]);
  assign or_1_cse = (fsm_output[2:1]!=2'b10);
  assign LOAD_DATA_OUTER_LOOP_len_not_4_nl = ~ z_out_1_32;
  assign LOAD_DATA_OUTER_LOOP_len_qr_6_0_lpi_2_dfm_1 = MUX_v_7_2_2(7'b0000000, (conf_info_crt_sva[6:0]),
      LOAD_DATA_OUTER_LOOP_len_not_4_nl);
  assign or_tmp_4 = (fsm_output[6:5]!=2'b00);
  assign and_tmp = (fsm_output[7]) & or_tmp_4;
  assign mux_tmp_2 = MUX_s_1_2_2(and_tmp, (fsm_output[7]), or_11_cse);
  assign mux_tmp_3 = MUX_s_1_2_2((~ or_tmp_4), or_tmp_4, fsm_output[7]);
  assign mux_tmp_4 = MUX_s_1_2_2(mux_tmp_3, (fsm_output[7]), or_11_cse);
  assign mux_tmp_5 = MUX_s_1_2_2(mux_tmp_4, mux_tmp_2, or_8_cse);
  assign mux_11_nl = MUX_s_1_2_2(mux_tmp_3, (fsm_output[7]), fsm_output[4]);
  assign mux_10_nl = MUX_s_1_2_2(and_tmp, (fsm_output[7]), fsm_output[4]);
  assign mux_tmp_8 = MUX_s_1_2_2(mux_11_nl, mux_10_nl, fsm_output[3]);
  assign and_dcpl_7 = (fsm_output[1:0]==2'b11);
  assign and_dcpl_8 = (fsm_output[3:2]==2'b01);
  assign and_dcpl_9 = and_dcpl_8 & and_dcpl_7;
  assign and_dcpl_10 = ~((fsm_output[7]) | (fsm_output[4]));
  assign and_dcpl_11 = (~ or_tmp_4) & and_dcpl_10;
  assign and_dcpl_13 = ~((fsm_output[1:0]!=2'b00));
  assign and_dcpl_14 = (fsm_output[3:2]==2'b10);
  assign and_dcpl_15 = and_dcpl_14 & and_dcpl_13;
  assign and_dcpl_17 = (fsm_output[1:0]==2'b01);
  assign and_dcpl_18 = and_dcpl_14 & and_dcpl_17;
  assign and_dcpl_20 = (fsm_output[1:0]==2'b10);
  assign and_dcpl_21 = and_dcpl_14 & and_dcpl_20;
  assign and_dcpl_23 = and_dcpl_14 & and_dcpl_7;
  assign and_dcpl_25 = (fsm_output[3:2]==2'b11);
  assign and_dcpl_26 = and_dcpl_25 & and_dcpl_13;
  assign and_dcpl_28 = and_dcpl_25 & and_dcpl_17;
  assign and_dcpl_30 = and_dcpl_25 & and_dcpl_20;
  assign and_dcpl_32 = and_dcpl_25 & and_dcpl_7;
  assign and_dcpl_34 = ~((fsm_output[3:2]!=2'b00));
  assign and_dcpl_35 = and_dcpl_34 & and_dcpl_13;
  assign and_dcpl_36 = (~ (fsm_output[7])) & (fsm_output[4]);
  assign and_dcpl_37 = (~ or_tmp_4) & and_dcpl_36;
  assign and_dcpl_39 = and_dcpl_34 & and_dcpl_17;
  assign and_dcpl_41 = and_dcpl_34 & and_dcpl_20;
  assign and_dcpl_43 = and_dcpl_34 & and_dcpl_7;
  assign and_dcpl_45 = and_dcpl_8 & and_dcpl_13;
  assign and_dcpl_47 = and_dcpl_8 & and_dcpl_17;
  assign and_dcpl_49 = and_dcpl_8 & and_dcpl_20;
  assign and_dcpl_60 = (fsm_output[6:5]==2'b01);
  assign and_dcpl_61 = and_dcpl_60 & and_dcpl_10;
  assign and_dcpl_78 = and_dcpl_60 & and_dcpl_36;
  assign and_dcpl_95 = (fsm_output[6:5]==2'b10);
  assign and_dcpl_96 = and_dcpl_95 & and_dcpl_10;
  assign and_dcpl_113 = and_dcpl_95 & and_dcpl_36;
  assign and_dcpl_130 = (fsm_output[6:5]==2'b11);
  assign and_dcpl_131 = and_dcpl_130 & and_dcpl_10;
  assign and_dcpl_148 = and_dcpl_130 & and_dcpl_36;
  assign and_dcpl_166 = (~ or_tmp_4) & (fsm_output[7]) & (~ (fsm_output[4]));
  assign and_dcpl_170 = and_dcpl_166 & and_dcpl_43;
  assign and_dcpl_175 = (fsm_output[2:0]==3'b101);
  assign and_dcpl_179 = (~ or_tmp_4) & (~ (fsm_output[7])) & nor_6_cse;
  assign or_dcpl_5 = (fsm_output[1:0]!=2'b10);
  assign or_dcpl_6 = (fsm_output[3:2]!=2'b01);
  assign or_dcpl_7 = or_dcpl_6 | or_dcpl_5;
  assign or_dcpl_9 = or_tmp_4 | (~ (fsm_output[7])) | (fsm_output[4]);
  assign and_dcpl_187 = and_dcpl_166 & and_dcpl_15;
  assign and_dcpl_188 = and_dcpl_11 & and_dcpl_39;
  assign and_dcpl_189 = and_dcpl_11 & and_dcpl_49;
  assign or_dcpl_21 = ~((fsm_output[1:0]==2'b11));
  assign or_dcpl_22 = (fsm_output[3:2]!=2'b00);
  assign or_dcpl_23 = or_dcpl_22 | or_dcpl_21;
  assign or_dcpl_24 = (fsm_output[7]) | (fsm_output[4]);
  assign or_dcpl_25 = or_tmp_4 | or_dcpl_24;
  assign and_dcpl_202 = and_dcpl_11 & and_dcpl_47;
  assign or_dcpl_32 = or_dcpl_6 | or_dcpl_21;
  assign or_dcpl_34 = (fsm_output[1:0]!=2'b00);
  assign or_dcpl_35 = (fsm_output[3:2]!=2'b10);
  assign or_dcpl_36 = or_dcpl_35 | or_dcpl_34;
  assign or_dcpl_38 = (fsm_output[1:0]!=2'b01);
  assign or_dcpl_39 = or_dcpl_35 | or_dcpl_38;
  assign or_dcpl_41 = or_dcpl_35 | or_dcpl_5;
  assign or_dcpl_43 = or_dcpl_35 | or_dcpl_21;
  assign or_dcpl_45 = ~((fsm_output[3:2]==2'b11));
  assign or_dcpl_46 = or_dcpl_45 | or_dcpl_34;
  assign or_dcpl_48 = or_dcpl_45 | or_dcpl_38;
  assign or_dcpl_50 = or_dcpl_45 | or_dcpl_5;
  assign or_dcpl_52 = or_dcpl_45 | or_dcpl_21;
  assign or_dcpl_54 = or_dcpl_22 | or_dcpl_34;
  assign or_dcpl_55 = (fsm_output[7]) | (~ (fsm_output[4]));
  assign or_dcpl_56 = or_tmp_4 | or_dcpl_55;
  assign or_dcpl_58 = or_dcpl_22 | or_dcpl_38;
  assign or_dcpl_60 = or_dcpl_22 | or_dcpl_5;
  assign or_dcpl_63 = or_dcpl_6 | or_dcpl_34;
  assign or_dcpl_65 = or_dcpl_6 | or_dcpl_38;
  assign or_dcpl_77 = (fsm_output[6:5]!=2'b01);
  assign or_dcpl_78 = or_dcpl_77 | or_dcpl_24;
  assign or_dcpl_95 = or_dcpl_77 | or_dcpl_55;
  assign or_dcpl_112 = (fsm_output[6:5]!=2'b10);
  assign or_dcpl_113 = or_dcpl_112 | or_dcpl_24;
  assign or_dcpl_130 = or_dcpl_112 | or_dcpl_55;
  assign or_dcpl_147 = ~((fsm_output[6:5]==2'b11));
  assign or_dcpl_148 = or_dcpl_147 | or_dcpl_24;
  assign or_dcpl_165 = or_dcpl_147 | or_dcpl_55;
  assign LOAD_DATA_INNER_LOOP_stage_0_mx0c0 = and_dcpl_11 & and_dcpl_45;
  assign LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_d_d = dma_read_chnl_Pop_mioi_return_rsc_z_mxwt;
  assign and_13_nl = and_dcpl_11 & and_dcpl_9;
  assign and_17_nl = and_dcpl_11 & and_dcpl_15;
  assign and_20_nl = and_dcpl_11 & and_dcpl_18;
  assign and_23_nl = and_dcpl_11 & and_dcpl_21;
  assign and_25_nl = and_dcpl_11 & and_dcpl_23;
  assign and_28_nl = and_dcpl_11 & and_dcpl_26;
  assign and_30_nl = and_dcpl_11 & and_dcpl_28;
  assign and_32_nl = and_dcpl_11 & and_dcpl_30;
  assign and_34_nl = and_dcpl_11 & and_dcpl_32;
  assign and_39_nl = and_dcpl_37 & and_dcpl_35;
  assign and_41_nl = and_dcpl_37 & and_dcpl_39;
  assign and_43_nl = and_dcpl_37 & and_dcpl_41;
  assign and_45_nl = and_dcpl_37 & and_dcpl_43;
  assign and_47_nl = and_dcpl_37 & and_dcpl_45;
  assign and_49_nl = and_dcpl_37 & and_dcpl_47;
  assign and_51_nl = and_dcpl_37 & and_dcpl_49;
  assign and_52_nl = and_dcpl_37 & and_dcpl_9;
  assign and_53_nl = and_dcpl_37 & and_dcpl_15;
  assign and_54_nl = and_dcpl_37 & and_dcpl_18;
  assign and_55_nl = and_dcpl_37 & and_dcpl_21;
  assign and_56_nl = and_dcpl_37 & and_dcpl_23;
  assign and_57_nl = and_dcpl_37 & and_dcpl_26;
  assign and_58_nl = and_dcpl_37 & and_dcpl_28;
  assign and_59_nl = and_dcpl_37 & and_dcpl_30;
  assign and_60_nl = and_dcpl_37 & and_dcpl_32;
  assign and_63_nl = and_dcpl_61 & and_dcpl_35;
  assign and_64_nl = and_dcpl_61 & and_dcpl_39;
  assign and_65_nl = and_dcpl_61 & and_dcpl_41;
  assign and_66_nl = and_dcpl_61 & and_dcpl_43;
  assign and_67_nl = and_dcpl_61 & and_dcpl_45;
  assign and_68_nl = and_dcpl_61 & and_dcpl_47;
  assign and_69_nl = and_dcpl_61 & and_dcpl_49;
  assign and_70_nl = and_dcpl_61 & and_dcpl_9;
  assign and_71_nl = and_dcpl_61 & and_dcpl_15;
  assign and_72_nl = and_dcpl_61 & and_dcpl_18;
  assign and_73_nl = and_dcpl_61 & and_dcpl_21;
  assign and_74_nl = and_dcpl_61 & and_dcpl_23;
  assign and_75_nl = and_dcpl_61 & and_dcpl_26;
  assign and_76_nl = and_dcpl_61 & and_dcpl_28;
  assign and_77_nl = and_dcpl_61 & and_dcpl_30;
  assign and_78_nl = and_dcpl_61 & and_dcpl_32;
  assign and_80_nl = and_dcpl_78 & and_dcpl_35;
  assign and_81_nl = and_dcpl_78 & and_dcpl_39;
  assign and_82_nl = and_dcpl_78 & and_dcpl_41;
  assign and_83_nl = and_dcpl_78 & and_dcpl_43;
  assign and_84_nl = and_dcpl_78 & and_dcpl_45;
  assign and_85_nl = and_dcpl_78 & and_dcpl_47;
  assign and_86_nl = and_dcpl_78 & and_dcpl_49;
  assign and_87_nl = and_dcpl_78 & and_dcpl_9;
  assign and_88_nl = and_dcpl_78 & and_dcpl_15;
  assign and_89_nl = and_dcpl_78 & and_dcpl_18;
  assign and_90_nl = and_dcpl_78 & and_dcpl_21;
  assign and_91_nl = and_dcpl_78 & and_dcpl_23;
  assign and_92_nl = and_dcpl_78 & and_dcpl_26;
  assign and_93_nl = and_dcpl_78 & and_dcpl_28;
  assign and_94_nl = and_dcpl_78 & and_dcpl_30;
  assign and_95_nl = and_dcpl_78 & and_dcpl_32;
  assign and_98_nl = and_dcpl_96 & and_dcpl_35;
  assign and_99_nl = and_dcpl_96 & and_dcpl_39;
  assign and_100_nl = and_dcpl_96 & and_dcpl_41;
  assign and_101_nl = and_dcpl_96 & and_dcpl_43;
  assign and_102_nl = and_dcpl_96 & and_dcpl_45;
  assign and_103_nl = and_dcpl_96 & and_dcpl_47;
  assign and_104_nl = and_dcpl_96 & and_dcpl_49;
  assign and_105_nl = and_dcpl_96 & and_dcpl_9;
  assign and_106_nl = and_dcpl_96 & and_dcpl_15;
  assign and_107_nl = and_dcpl_96 & and_dcpl_18;
  assign and_108_nl = and_dcpl_96 & and_dcpl_21;
  assign and_109_nl = and_dcpl_96 & and_dcpl_23;
  assign and_110_nl = and_dcpl_96 & and_dcpl_26;
  assign and_111_nl = and_dcpl_96 & and_dcpl_28;
  assign and_112_nl = and_dcpl_96 & and_dcpl_30;
  assign and_113_nl = and_dcpl_96 & and_dcpl_32;
  assign and_115_nl = and_dcpl_113 & and_dcpl_35;
  assign and_116_nl = and_dcpl_113 & and_dcpl_39;
  assign and_117_nl = and_dcpl_113 & and_dcpl_41;
  assign and_118_nl = and_dcpl_113 & and_dcpl_43;
  assign and_119_nl = and_dcpl_113 & and_dcpl_45;
  assign and_120_nl = and_dcpl_113 & and_dcpl_47;
  assign and_121_nl = and_dcpl_113 & and_dcpl_49;
  assign and_122_nl = and_dcpl_113 & and_dcpl_9;
  assign and_123_nl = and_dcpl_113 & and_dcpl_15;
  assign and_124_nl = and_dcpl_113 & and_dcpl_18;
  assign and_125_nl = and_dcpl_113 & and_dcpl_21;
  assign and_126_nl = and_dcpl_113 & and_dcpl_23;
  assign and_127_nl = and_dcpl_113 & and_dcpl_26;
  assign and_128_nl = and_dcpl_113 & and_dcpl_28;
  assign and_129_nl = and_dcpl_113 & and_dcpl_30;
  assign and_130_nl = and_dcpl_113 & and_dcpl_32;
  assign and_133_nl = and_dcpl_131 & and_dcpl_35;
  assign and_134_nl = and_dcpl_131 & and_dcpl_39;
  assign and_135_nl = and_dcpl_131 & and_dcpl_41;
  assign and_136_nl = and_dcpl_131 & and_dcpl_43;
  assign and_137_nl = and_dcpl_131 & and_dcpl_45;
  assign and_138_nl = and_dcpl_131 & and_dcpl_47;
  assign and_139_nl = and_dcpl_131 & and_dcpl_49;
  assign and_140_nl = and_dcpl_131 & and_dcpl_9;
  assign and_141_nl = and_dcpl_131 & and_dcpl_15;
  assign and_142_nl = and_dcpl_131 & and_dcpl_18;
  assign and_143_nl = and_dcpl_131 & and_dcpl_21;
  assign and_144_nl = and_dcpl_131 & and_dcpl_23;
  assign and_145_nl = and_dcpl_131 & and_dcpl_26;
  assign and_146_nl = and_dcpl_131 & and_dcpl_28;
  assign and_147_nl = and_dcpl_131 & and_dcpl_30;
  assign and_148_nl = and_dcpl_131 & and_dcpl_32;
  assign and_150_nl = and_dcpl_148 & and_dcpl_35;
  assign and_151_nl = and_dcpl_148 & and_dcpl_39;
  assign and_152_nl = and_dcpl_148 & and_dcpl_41;
  assign and_153_nl = and_dcpl_148 & and_dcpl_43;
  assign and_154_nl = and_dcpl_148 & and_dcpl_45;
  assign and_155_nl = and_dcpl_148 & and_dcpl_47;
  assign and_156_nl = and_dcpl_148 & and_dcpl_49;
  assign and_157_nl = and_dcpl_148 & and_dcpl_9;
  assign and_158_nl = and_dcpl_148 & and_dcpl_15;
  assign and_159_nl = and_dcpl_148 & and_dcpl_18;
  assign and_160_nl = and_dcpl_148 & and_dcpl_21;
  assign and_161_nl = and_dcpl_148 & and_dcpl_23;
  assign and_162_nl = and_dcpl_148 & and_dcpl_26;
  assign and_163_nl = and_dcpl_148 & and_dcpl_28;
  assign and_164_nl = and_dcpl_148 & and_dcpl_30;
  assign and_165_nl = and_dcpl_148 & and_dcpl_32;
  assign and_168_nl = and_dcpl_166 & and_dcpl_35;
  assign and_169_nl = and_dcpl_166 & and_dcpl_39;
  assign and_170_nl = and_dcpl_166 & and_dcpl_41;
  assign and_172_nl = and_dcpl_166 & and_dcpl_45;
  assign mux1h_nl = MUX1HOT_v_7_126_2(7'b1111110, 7'b1111101, 7'b1111100, 7'b1111011,
      7'b1111010, 7'b1111001, 7'b1111000, 7'b1110111, 7'b1110110, 7'b1110101, 7'b1110100,
      7'b1110011, 7'b1110010, 7'b1110001, 7'b1110000, 7'b1101111, 7'b1101110, 7'b1101101,
      7'b1101100, 7'b1101011, 7'b1101010, 7'b1101001, 7'b1101000, 7'b1100111, 7'b1100110,
      7'b1100101, 7'b1100100, 7'b1100011, 7'b1100010, 7'b1100001, 7'b1100000, 7'b1011111,
      7'b1011110, 7'b1011101, 7'b1011100, 7'b1011011, 7'b1011010, 7'b1011001, 7'b1011000,
      7'b1010111, 7'b1010110, 7'b1010101, 7'b1010100, 7'b1010011, 7'b1010010, 7'b1010001,
      7'b1010000, 7'b1001111, 7'b1001110, 7'b1001101, 7'b1001100, 7'b1001011, 7'b1001010,
      7'b1001001, 7'b1001000, 7'b1000111, 7'b1000110, 7'b1000101, 7'b1000100, 7'b1000011,
      7'b1000010, 7'b1000001, 7'b1000000, 7'b0111111, 7'b0111110, 7'b0111101, 7'b0111100,
      7'b0111011, 7'b0111010, 7'b0111001, 7'b0111000, 7'b0110111, 7'b0110110, 7'b0110101,
      7'b0110100, 7'b0110011, 7'b0110010, 7'b0110001, 7'b0110000, 7'b0101111, 7'b0101110,
      7'b0101101, 7'b0101100, 7'b0101011, 7'b0101010, 7'b0101001, 7'b0101000, 7'b0100111,
      7'b0100110, 7'b0100101, 7'b0100100, 7'b0100011, 7'b0100010, 7'b0100001, 7'b0100000,
      7'b0011111, 7'b0011110, 7'b0011101, 7'b0011100, 7'b0011011, 7'b0011010, 7'b0011001,
      7'b0011000, 7'b0010111, 7'b0010110, 7'b0010101, 7'b0010100, 7'b0010011, 7'b0010010,
      7'b0010001, 7'b0010000, 7'b0001111, 7'b0001110, 7'b0001101, 7'b0001100, 7'b0001011,
      7'b0001010, 7'b0001001, 7'b0001000, 7'b0000111, 7'b0000110, 7'b0000101, 7'b0000100,
      7'b0000011, 7'b0000010, 7'b0000001, {and_13_nl , and_17_nl , and_20_nl , and_23_nl
      , and_25_nl , and_28_nl , and_30_nl , and_32_nl , and_34_nl , and_39_nl , and_41_nl
      , and_43_nl , and_45_nl , and_47_nl , and_49_nl , and_51_nl , and_52_nl , and_53_nl
      , and_54_nl , and_55_nl , and_56_nl , and_57_nl , and_58_nl , and_59_nl , and_60_nl
      , and_63_nl , and_64_nl , and_65_nl , and_66_nl , and_67_nl , and_68_nl , and_69_nl
      , and_70_nl , and_71_nl , and_72_nl , and_73_nl , and_74_nl , and_75_nl , and_76_nl
      , and_77_nl , and_78_nl , and_80_nl , and_81_nl , and_82_nl , and_83_nl , and_84_nl
      , and_85_nl , and_86_nl , and_87_nl , and_88_nl , and_89_nl , and_90_nl , and_91_nl
      , and_92_nl , and_93_nl , and_94_nl , and_95_nl , and_98_nl , and_99_nl , and_100_nl
      , and_101_nl , and_102_nl , and_103_nl , and_104_nl , and_105_nl , and_106_nl
      , and_107_nl , and_108_nl , and_109_nl , and_110_nl , and_111_nl , and_112_nl
      , and_113_nl , and_115_nl , and_116_nl , and_117_nl , and_118_nl , and_119_nl
      , and_120_nl , and_121_nl , and_122_nl , and_123_nl , and_124_nl , and_125_nl
      , and_126_nl , and_127_nl , and_128_nl , and_129_nl , and_130_nl , and_133_nl
      , and_134_nl , and_135_nl , and_136_nl , and_137_nl , and_138_nl , and_139_nl
      , and_140_nl , and_141_nl , and_142_nl , and_143_nl , and_144_nl , and_145_nl
      , and_146_nl , and_147_nl , and_148_nl , and_150_nl , and_151_nl , and_152_nl
      , and_153_nl , and_154_nl , and_155_nl , and_156_nl , and_157_nl , and_158_nl
      , and_159_nl , and_160_nl , and_161_nl , and_162_nl , and_163_nl , and_164_nl
      , and_165_nl , and_168_nl , and_169_nl , and_170_nl , and_dcpl_170 , and_172_nl});
  assign or_12_nl = (fsm_output[7]) | (~ or_tmp_4);
  assign mux_25_nl = MUX_s_1_2_2(or_12_nl, (fsm_output[7]), or_11_cse);
  assign mux_27_nl = MUX_s_1_2_2(mux_tmp_4, mux_25_nl, and_205_cse);
  assign or_9_nl = and_205_cse | (fsm_output[4:3]!=2'b00);
  assign mux_24_nl = MUX_s_1_2_2(mux_tmp_3, (fsm_output[7]), or_9_nl);
  assign mux_28_nl = MUX_s_1_2_2(mux_27_nl, mux_24_nl, fsm_output[0]);
  assign nor_12_nl = ~(MUX_v_7_2_2(mux1h_nl, 7'b1111111, mux_28_nl));
  assign and_173_nl = and_dcpl_166 & and_dcpl_47;
  assign LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_radr_d = MUX_v_7_2_2(nor_12_nl,
      7'b1111111, and_173_nl);
  assign LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_wadr_d = LOAD_DATA_INNER_LOOP_slc_LOAD_DATA_INNER_LOOP_i_6_0_itm_1;
  assign LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_we_d_pff = and_dcpl_179 & and_dcpl_175
      & LOAD_DATA_INNER_LOOP_stage_0_2 & (~ exit_LOAD_DATA_INNER_LOOP_sva_st_1);
  assign LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = (or_tmp_4 | (fsm_output[4]) | and_205_cse | (fsm_output[3])) ^ (fsm_output[7]);
  assign nor_16_cse = ~((fsm_output[6:5]!=2'b00));
  assign and_dcpl_214 = (fsm_output[4:3]==2'b01) & nor_16_cse & (fsm_output[7]) &
      (~ (fsm_output[1])) & (~ (fsm_output[2])) & (~ (fsm_output[0]));
  assign and_dcpl_215 = (~ (fsm_output[2])) & (fsm_output[0]);
  assign and_dcpl_216 = ~((fsm_output[7]) | (fsm_output[1]));
  assign and_dcpl_219 = ~((fsm_output[4]) | (fsm_output[6]));
  assign and_dcpl_220 = and_dcpl_219 & (~ (fsm_output[5])) & (~ (fsm_output[3]));
  assign and_dcpl_221 = and_dcpl_220 & and_dcpl_216 & and_dcpl_215;
  assign and_dcpl_222 = ~((fsm_output[2]) | (fsm_output[0]));
  assign and_dcpl_227 = and_dcpl_219 & (~ (fsm_output[5])) & (fsm_output[3]) & (fsm_output[7])
      & (~ (fsm_output[1])) & and_dcpl_222;
  assign and_dcpl_228 = (~ (fsm_output[7])) & (fsm_output[1]);
  assign and_dcpl_230 = and_dcpl_220 & and_dcpl_228 & and_dcpl_215;
  assign and_dcpl_233 = and_dcpl_220 & and_dcpl_216 & (fsm_output[2]) & (fsm_output[0]);
  assign and_dcpl_235 = and_dcpl_220 & and_dcpl_228 & and_dcpl_222;
  assign and_dcpl_238 = and_dcpl_220 & and_dcpl_228 & (fsm_output[2]) & (~ (fsm_output[0]));
  assign and_dcpl_249 = nor_6_cse & nor_16_cse & (~ (fsm_output[7])) & (fsm_output[1])
      & (fsm_output[2]) & (~ (fsm_output[0]));
  assign LOAD_BATCH_LOOP_or_1_ssc = and_dcpl_221 | and_dcpl_235 | and_dcpl_238;
  always @(posedge clk) begin
    if ( load_input_wen ) begin
      conf_info_crt_sva <= MUX_v_64_2_2(conf_info_crt_sva, conf_info, mux_35_nl);
      offset_lpi_2 <= MUX_v_32_2_2(32'b00000000000000000000000000000000, LOAD_BATCH_LOOP_b_mux_nl,
          not_nl);
      LOAD_DATA_OUTER_LOOP_s_31_7_sva <= MUX1HOT_v_25_3_2((conf_info_crt_sva[31:7]),
          z_out_2, LOAD_DATA_OUTER_LOOP_s_31_7_sva, {and_192_nl , and_dcpl_189 ,
          (~ mux_42_nl)});
      LOAD_DATA_INNER_LOOP_i_sva <= MUX_v_16_2_2(16'b0000000000000000, (z_out_2[15:0]),
          and_dcpl_202);
      LOAD_DATA_INNER_LOOP_slc_LOAD_DATA_INNER_LOOP_i_6_0_itm_1 <= LOAD_DATA_INNER_LOOP_i_sva[6:0];
      LOAD_DATA_OUTER_LOOP_asn_8_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      reg_dma_read_ctrl_Push_mioi_oswt_cse <= 1'b0;
      reg_dma_read_chnl_Pop_mioi_oswt_cse <= 1'b0;
      reg_input_ready_channel_Pop_mioi_oswt_cse <= 1'b0;
      exit_LOAD_DATA_INNER_LOOP_sva_st_1 <= 1'b0;
      LOAD_DATA_INNER_LOOP_stage_0_2 <= 1'b0;
    end
    else if ( load_input_wen ) begin
      reg_dma_read_ctrl_Push_mioi_oswt_cse <= and_183_rmff;
      reg_dma_read_chnl_Pop_mioi_oswt_cse <= and_186_rmff;
      reg_input_ready_channel_Pop_mioi_oswt_cse <= and_187_rmff;
      exit_LOAD_DATA_INNER_LOOP_sva_st_1 <= ~ z_out_1_32;
      LOAD_DATA_INNER_LOOP_stage_0_2 <= LOAD_DATA_INNER_LOOP_stage_0 & and_dcpl_202;
    end
  end
  always @(posedge clk) begin
    if ( LOAD_DATA_OUTER_LOOP_and_cse ) begin
      plm_in_cnsi_idat_2047_2016 <= LOAD_DATA_OUTER_LOOP_asn_71_itm;
      plm_in_cnsi_idat_2079_2048 <= LOAD_DATA_OUTER_LOOP_asn_70_itm;
      plm_in_cnsi_idat_2015_1984 <= LOAD_DATA_OUTER_LOOP_asn_72_itm;
      plm_in_cnsi_idat_2111_2080 <= LOAD_DATA_OUTER_LOOP_asn_69_itm;
      plm_in_cnsi_idat_1983_1952 <= LOAD_DATA_OUTER_LOOP_asn_73_itm;
      plm_in_cnsi_idat_2143_2112 <= LOAD_DATA_OUTER_LOOP_asn_68_itm;
      plm_in_cnsi_idat_1951_1920 <= LOAD_DATA_OUTER_LOOP_asn_74_itm;
      plm_in_cnsi_idat_2175_2144 <= LOAD_DATA_OUTER_LOOP_asn_67_itm;
      plm_in_cnsi_idat_1919_1888 <= LOAD_DATA_OUTER_LOOP_asn_75_itm;
      plm_in_cnsi_idat_2207_2176 <= LOAD_DATA_OUTER_LOOP_asn_66_itm;
      plm_in_cnsi_idat_1887_1856 <= LOAD_DATA_OUTER_LOOP_asn_76_itm;
      plm_in_cnsi_idat_2239_2208 <= LOAD_DATA_OUTER_LOOP_asn_65_itm;
      plm_in_cnsi_idat_1855_1824 <= LOAD_DATA_OUTER_LOOP_asn_77_itm;
      plm_in_cnsi_idat_2271_2240 <= LOAD_DATA_OUTER_LOOP_asn_64_itm;
      plm_in_cnsi_idat_1823_1792 <= LOAD_DATA_OUTER_LOOP_asn_78_itm;
      plm_in_cnsi_idat_2303_2272 <= LOAD_DATA_OUTER_LOOP_asn_63_itm;
      plm_in_cnsi_idat_1791_1760 <= LOAD_DATA_OUTER_LOOP_asn_79_itm;
      plm_in_cnsi_idat_2335_2304 <= LOAD_DATA_OUTER_LOOP_asn_62_itm;
      plm_in_cnsi_idat_1759_1728 <= LOAD_DATA_OUTER_LOOP_asn_80_itm;
      plm_in_cnsi_idat_2367_2336 <= LOAD_DATA_OUTER_LOOP_asn_61_itm;
      plm_in_cnsi_idat_1727_1696 <= LOAD_DATA_OUTER_LOOP_asn_81_itm;
      plm_in_cnsi_idat_2399_2368 <= LOAD_DATA_OUTER_LOOP_asn_60_itm;
      plm_in_cnsi_idat_1695_1664 <= LOAD_DATA_OUTER_LOOP_asn_82_itm;
      plm_in_cnsi_idat_2431_2400 <= LOAD_DATA_OUTER_LOOP_asn_59_itm;
      plm_in_cnsi_idat_1663_1632 <= LOAD_DATA_OUTER_LOOP_asn_83_itm;
      plm_in_cnsi_idat_2463_2432 <= LOAD_DATA_OUTER_LOOP_asn_58_itm;
      plm_in_cnsi_idat_1631_1600 <= LOAD_DATA_OUTER_LOOP_asn_84_itm;
      plm_in_cnsi_idat_2495_2464 <= LOAD_DATA_OUTER_LOOP_asn_57_itm;
      plm_in_cnsi_idat_1599_1568 <= LOAD_DATA_OUTER_LOOP_asn_85_itm;
      plm_in_cnsi_idat_2527_2496 <= LOAD_DATA_OUTER_LOOP_asn_56_itm;
      plm_in_cnsi_idat_1567_1536 <= LOAD_DATA_OUTER_LOOP_asn_86_itm;
      plm_in_cnsi_idat_2559_2528 <= LOAD_DATA_OUTER_LOOP_asn_55_itm;
      plm_in_cnsi_idat_1535_1504 <= LOAD_DATA_OUTER_LOOP_asn_87_itm;
      plm_in_cnsi_idat_2591_2560 <= LOAD_DATA_OUTER_LOOP_asn_54_itm;
      plm_in_cnsi_idat_1503_1472 <= LOAD_DATA_OUTER_LOOP_asn_88_itm;
      plm_in_cnsi_idat_2623_2592 <= LOAD_DATA_OUTER_LOOP_asn_53_itm;
      plm_in_cnsi_idat_1471_1440 <= LOAD_DATA_OUTER_LOOP_asn_89_itm;
      plm_in_cnsi_idat_2655_2624 <= LOAD_DATA_OUTER_LOOP_asn_52_itm;
      plm_in_cnsi_idat_1439_1408 <= LOAD_DATA_OUTER_LOOP_asn_90_itm;
      plm_in_cnsi_idat_2687_2656 <= LOAD_DATA_OUTER_LOOP_asn_51_itm;
      plm_in_cnsi_idat_1407_1376 <= LOAD_DATA_OUTER_LOOP_asn_91_itm;
      plm_in_cnsi_idat_2719_2688 <= LOAD_DATA_OUTER_LOOP_asn_50_itm;
      plm_in_cnsi_idat_1375_1344 <= LOAD_DATA_OUTER_LOOP_asn_92_itm;
      plm_in_cnsi_idat_2751_2720 <= LOAD_DATA_OUTER_LOOP_asn_49_itm;
      plm_in_cnsi_idat_1343_1312 <= LOAD_DATA_OUTER_LOOP_asn_93_itm;
      plm_in_cnsi_idat_2783_2752 <= LOAD_DATA_OUTER_LOOP_asn_48_itm;
      plm_in_cnsi_idat_1311_1280 <= LOAD_DATA_OUTER_LOOP_asn_94_itm;
      plm_in_cnsi_idat_2815_2784 <= LOAD_DATA_OUTER_LOOP_asn_47_itm;
      plm_in_cnsi_idat_1279_1248 <= LOAD_DATA_OUTER_LOOP_asn_95_itm;
      plm_in_cnsi_idat_2847_2816 <= LOAD_DATA_OUTER_LOOP_asn_46_itm;
      plm_in_cnsi_idat_1247_1216 <= LOAD_DATA_OUTER_LOOP_asn_96_itm;
      plm_in_cnsi_idat_2879_2848 <= LOAD_DATA_OUTER_LOOP_asn_45_itm;
      plm_in_cnsi_idat_1215_1184 <= LOAD_DATA_OUTER_LOOP_asn_97_itm;
      plm_in_cnsi_idat_2911_2880 <= LOAD_DATA_OUTER_LOOP_asn_44_itm;
      plm_in_cnsi_idat_1183_1152 <= LOAD_DATA_OUTER_LOOP_asn_98_itm;
      plm_in_cnsi_idat_2943_2912 <= LOAD_DATA_OUTER_LOOP_asn_43_itm;
      plm_in_cnsi_idat_1151_1120 <= LOAD_DATA_OUTER_LOOP_asn_99_itm;
      plm_in_cnsi_idat_2975_2944 <= LOAD_DATA_OUTER_LOOP_asn_42_itm;
      plm_in_cnsi_idat_1119_1088 <= LOAD_DATA_OUTER_LOOP_asn_100_itm;
      plm_in_cnsi_idat_3007_2976 <= LOAD_DATA_OUTER_LOOP_asn_41_itm;
      plm_in_cnsi_idat_1087_1056 <= LOAD_DATA_OUTER_LOOP_asn_101_itm;
      plm_in_cnsi_idat_3039_3008 <= LOAD_DATA_OUTER_LOOP_asn_40_itm;
      plm_in_cnsi_idat_1055_1024 <= LOAD_DATA_OUTER_LOOP_asn_102_itm;
      plm_in_cnsi_idat_3071_3040 <= LOAD_DATA_OUTER_LOOP_asn_39_itm;
      plm_in_cnsi_idat_1023_992 <= LOAD_DATA_OUTER_LOOP_asn_103_itm;
      plm_in_cnsi_idat_3103_3072 <= LOAD_DATA_OUTER_LOOP_asn_38_itm;
      plm_in_cnsi_idat_991_960 <= LOAD_DATA_OUTER_LOOP_asn_104_itm;
      plm_in_cnsi_idat_3135_3104 <= LOAD_DATA_OUTER_LOOP_asn_37_itm;
      plm_in_cnsi_idat_959_928 <= LOAD_DATA_OUTER_LOOP_asn_105_itm;
      plm_in_cnsi_idat_3167_3136 <= LOAD_DATA_OUTER_LOOP_asn_36_itm;
      plm_in_cnsi_idat_927_896 <= LOAD_DATA_OUTER_LOOP_asn_106_itm;
      plm_in_cnsi_idat_3199_3168 <= LOAD_DATA_OUTER_LOOP_asn_35_itm;
      plm_in_cnsi_idat_895_864 <= LOAD_DATA_OUTER_LOOP_asn_107_itm;
      plm_in_cnsi_idat_3231_3200 <= LOAD_DATA_OUTER_LOOP_asn_34_itm;
      plm_in_cnsi_idat_863_832 <= LOAD_DATA_OUTER_LOOP_asn_108_itm;
      plm_in_cnsi_idat_3263_3232 <= LOAD_DATA_OUTER_LOOP_asn_33_itm;
      plm_in_cnsi_idat_831_800 <= LOAD_DATA_OUTER_LOOP_asn_109_itm;
      plm_in_cnsi_idat_3295_3264 <= LOAD_DATA_OUTER_LOOP_asn_32_itm;
      plm_in_cnsi_idat_799_768 <= LOAD_DATA_OUTER_LOOP_asn_110_itm;
      plm_in_cnsi_idat_3327_3296 <= LOAD_DATA_OUTER_LOOP_asn_31_itm;
      plm_in_cnsi_idat_767_736 <= LOAD_DATA_OUTER_LOOP_asn_111_itm;
      plm_in_cnsi_idat_3359_3328 <= LOAD_DATA_OUTER_LOOP_asn_30_itm;
      plm_in_cnsi_idat_735_704 <= LOAD_DATA_OUTER_LOOP_asn_112_itm;
      plm_in_cnsi_idat_3391_3360 <= LOAD_DATA_OUTER_LOOP_asn_29_itm;
      plm_in_cnsi_idat_703_672 <= LOAD_DATA_OUTER_LOOP_asn_113_itm;
      plm_in_cnsi_idat_3423_3392 <= LOAD_DATA_OUTER_LOOP_asn_28_itm;
      plm_in_cnsi_idat_671_640 <= LOAD_DATA_OUTER_LOOP_asn_114_itm;
      plm_in_cnsi_idat_3455_3424 <= LOAD_DATA_OUTER_LOOP_asn_27_itm;
      plm_in_cnsi_idat_639_608 <= LOAD_DATA_OUTER_LOOP_asn_115_itm;
      plm_in_cnsi_idat_3487_3456 <= LOAD_DATA_OUTER_LOOP_asn_26_itm;
      plm_in_cnsi_idat_607_576 <= LOAD_DATA_OUTER_LOOP_asn_116_itm;
      plm_in_cnsi_idat_3519_3488 <= LOAD_DATA_OUTER_LOOP_asn_25_itm;
      plm_in_cnsi_idat_575_544 <= LOAD_DATA_OUTER_LOOP_asn_117_itm;
      plm_in_cnsi_idat_3551_3520 <= LOAD_DATA_OUTER_LOOP_asn_24_itm;
      plm_in_cnsi_idat_543_512 <= LOAD_DATA_OUTER_LOOP_asn_118_itm;
      plm_in_cnsi_idat_3583_3552 <= LOAD_DATA_OUTER_LOOP_asn_23_itm;
      plm_in_cnsi_idat_511_480 <= LOAD_DATA_OUTER_LOOP_asn_119_itm;
      plm_in_cnsi_idat_3615_3584 <= LOAD_DATA_OUTER_LOOP_asn_22_itm;
      plm_in_cnsi_idat_479_448 <= LOAD_DATA_OUTER_LOOP_asn_120_itm;
      plm_in_cnsi_idat_3647_3616 <= LOAD_DATA_OUTER_LOOP_asn_21_itm;
      plm_in_cnsi_idat_447_416 <= LOAD_DATA_OUTER_LOOP_asn_121_itm;
      plm_in_cnsi_idat_3679_3648 <= LOAD_DATA_OUTER_LOOP_asn_20_itm;
      plm_in_cnsi_idat_415_384 <= LOAD_DATA_OUTER_LOOP_asn_122_itm;
      plm_in_cnsi_idat_3711_3680 <= LOAD_DATA_OUTER_LOOP_asn_19_itm;
      plm_in_cnsi_idat_383_352 <= LOAD_DATA_OUTER_LOOP_asn_123_itm;
      plm_in_cnsi_idat_3743_3712 <= LOAD_DATA_OUTER_LOOP_asn_18_itm;
      plm_in_cnsi_idat_351_320 <= LOAD_DATA_OUTER_LOOP_asn_124_itm;
      plm_in_cnsi_idat_3775_3744 <= LOAD_DATA_OUTER_LOOP_asn_17_itm;
      plm_in_cnsi_idat_319_288 <= LOAD_DATA_OUTER_LOOP_asn_125_itm;
      plm_in_cnsi_idat_3807_3776 <= LOAD_DATA_OUTER_LOOP_asn_16_itm;
      plm_in_cnsi_idat_287_256 <= LOAD_DATA_OUTER_LOOP_asn_126_itm;
      plm_in_cnsi_idat_3839_3808 <= LOAD_DATA_OUTER_LOOP_asn_15_itm;
      plm_in_cnsi_idat_255_224 <= LOAD_DATA_OUTER_LOOP_asn_127_itm;
      plm_in_cnsi_idat_3871_3840 <= LOAD_DATA_OUTER_LOOP_asn_14_itm;
      plm_in_cnsi_idat_223_192 <= LOAD_DATA_OUTER_LOOP_asn_128_itm;
      plm_in_cnsi_idat_3903_3872 <= LOAD_DATA_OUTER_LOOP_asn_13_itm;
      plm_in_cnsi_idat_191_160 <= LOAD_DATA_OUTER_LOOP_asn_129_itm;
      plm_in_cnsi_idat_3935_3904 <= LOAD_DATA_OUTER_LOOP_asn_12_itm;
      plm_in_cnsi_idat_159_128 <= LOAD_DATA_OUTER_LOOP_asn_130_itm;
      plm_in_cnsi_idat_3967_3936 <= LOAD_DATA_OUTER_LOOP_asn_11_itm;
      plm_in_cnsi_idat_127_96 <= LOAD_DATA_OUTER_LOOP_asn_131_itm;
      plm_in_cnsi_idat_3999_3968 <= LOAD_DATA_OUTER_LOOP_asn_10_itm;
      plm_in_cnsi_idat_95_64 <= LOAD_DATA_OUTER_LOOP_asn_132_itm;
      plm_in_cnsi_idat_4031_4000 <= LOAD_DATA_OUTER_LOOP_asn_9_itm;
      plm_in_cnsi_idat_63_32 <= LOAD_DATA_OUTER_LOOP_asn_133_itm;
      plm_in_cnsi_idat_4063_4032 <= LOAD_DATA_OUTER_LOOP_asn_8_itm;
      plm_in_cnsi_idat_31_0 <= LOAD_DATA_OUTER_LOOP_asn_134_itm;
      plm_in_cnsi_idat_4095_4064 <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (and_dcpl_188 | and_dcpl_187) ) begin
      LOAD_BATCH_LOOP_b_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000,
          z_out, and_dcpl_187);
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_25 | or_dcpl_23)) ) begin
      LOAD_DATA_OUTER_LOOP_len_qr_6_0_lpi_2_dfm <= LOAD_DATA_OUTER_LOOP_len_qr_6_0_lpi_2_dfm_1;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & ((~(mux_5_nl | (fsm_output[7:5]!=3'b000) | (~ nor_6_cse)))
        | and_dcpl_170) ) begin
      LOAD_DATA_OUTER_LOOP_asn_10_itm <= MUX_v_32_2_2(({7'b0000000 , LOAD_DATA_OUTER_LOOP_len_qif_mux1h_nl}),
          LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d, and_dcpl_170);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_DATA_INNER_LOOP_stage_0 <= 1'b0;
    end
    else if ( load_input_wen & (LOAD_DATA_INNER_LOOP_stage_0_mx0c0 | and_dcpl_202
        | and_dcpl_189) ) begin
      LOAD_DATA_INNER_LOOP_stage_0 <= LOAD_DATA_OUTER_LOOP_mux_nl | LOAD_DATA_INNER_LOOP_stage_0_mx0c0;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_25 | or_dcpl_32)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_134_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_25 | or_dcpl_36)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_133_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_25 | or_dcpl_39)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_132_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_25 | or_dcpl_41)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_131_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_25 | or_dcpl_43)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_130_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_25 | or_dcpl_46)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_129_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_25 | or_dcpl_48)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_128_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_25 | or_dcpl_50)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_127_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_25 | or_dcpl_52)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_126_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_54)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_125_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_58)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_124_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_60)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_123_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_23)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_122_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_63)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_121_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_65)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_120_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_7)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_119_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_32)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_118_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_36)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_117_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_39)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_116_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_41)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_115_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_43)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_114_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_46)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_113_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_48)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_112_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_50)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_111_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_56 | or_dcpl_52)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_110_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_54)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_109_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_58)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_108_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_60)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_107_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_23)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_106_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_63)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_105_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_65)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_104_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_7)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_103_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_32)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_102_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_36)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_101_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_39)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_100_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_41)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_99_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_43)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_98_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_46)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_97_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_48)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_96_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_50)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_95_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_78 | or_dcpl_52)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_94_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_54)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_93_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_58)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_92_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_60)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_91_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_23)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_90_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_63)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_89_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_65)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_88_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_7)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_87_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_32)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_86_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_36)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_85_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_39)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_84_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_41)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_83_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_43)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_82_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_46)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_81_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_48)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_80_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_50)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_79_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_95 | or_dcpl_52)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_78_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_54)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_77_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_58)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_76_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_60)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_75_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_23)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_74_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_63)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_73_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_65)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_72_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_7)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_71_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_32)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_70_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_36)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_69_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_39)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_68_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_41)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_67_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_43)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_66_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_46)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_65_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_48)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_64_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_50)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_63_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_113 | or_dcpl_52)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_62_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_54)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_61_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_58)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_60_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_60)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_59_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_23)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_58_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_63)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_57_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_65)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_56_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_7)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_55_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_32)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_54_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_36)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_53_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_39)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_52_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_41)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_51_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_43)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_50_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_46)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_49_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_48)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_48_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_50)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_47_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_130 | or_dcpl_52)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_46_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_54)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_45_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_58)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_44_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_60)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_43_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_23)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_42_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_63)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_41_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_65)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_40_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_7)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_39_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_32)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_38_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_36)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_37_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_39)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_36_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_41)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_35_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_43)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_34_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_46)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_33_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_48)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_32_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_50)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_31_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_148 | or_dcpl_52)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_30_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_54)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_29_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_58)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_28_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_60)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_27_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_23)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_26_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_63)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_25_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_65)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_24_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_7)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_23_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_32)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_22_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_36)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_21_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_39)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_20_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_41)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_19_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_43)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_18_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_46)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_17_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_48)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_16_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_50)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_15_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_165 | or_dcpl_52)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_14_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_9 | or_dcpl_54)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_13_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_9 | or_dcpl_58)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_12_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_9 | or_dcpl_60)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_11_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( load_input_wen & (~(or_dcpl_9 | or_dcpl_63)) ) begin
      LOAD_DATA_OUTER_LOOP_asn_9_itm <= LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
    end
  end
  assign mux_13_nl = MUX_s_1_2_2(mux_tmp_8, mux_tmp_2, or_8_cse);
  assign mux_35_nl = MUX_s_1_2_2(mux_13_nl, mux_tmp_5, fsm_output[0]);
  assign mux_19_nl = MUX_s_1_2_2(mux_tmp_8, mux_tmp_2, fsm_output[2]);
  assign mux_37_nl = MUX_s_1_2_2(mux_tmp_2, mux_tmp_4, fsm_output[2]);
  assign mux_20_nl = MUX_s_1_2_2(mux_19_nl, mux_37_nl, fsm_output[1]);
  assign mux_21_nl = MUX_s_1_2_2(mux_20_nl, mux_tmp_5, fsm_output[0]);
  assign LOAD_BATCH_LOOP_b_mux_nl = MUX_v_32_2_2(offset_lpi_2, z_out, mux_21_nl);
  assign not_nl = ~ and_dcpl_188;
  assign and_192_nl = and_dcpl_11 & and_dcpl_41;
  assign nor_3_nl = ~((fsm_output[2:1]!=2'b10));
  assign mux_41_nl = MUX_s_1_2_2(mux_tmp_4, mux_tmp_2, nor_3_nl);
  assign mux_42_nl = MUX_s_1_2_2(mux_41_nl, mux_tmp_5, fsm_output[0]);
  assign nor_4_nl = ~(z_out_1_32 | (~ (fsm_output[0])));
  assign mux_44_nl = MUX_s_1_2_2(or_1_cse, mux_4_cse, nor_4_nl);
  assign or_37_nl = mux_44_nl | (fsm_output[7:5]!=3'b000) | or_11_cse;
  assign and_196_nl = and_dcpl_179 & (fsm_output[2:0]==3'b011) & (~ z_out_1_32);
  assign and_198_nl = and_dcpl_11 & and_dcpl_8 & (~ (fsm_output[1]));
  assign LOAD_DATA_OUTER_LOOP_len_qif_mux1h_nl = MUX1HOT_v_25_3_2(25'b0000000000000000000000001,
      LOAD_DATA_OUTER_LOOP_s_31_7_sva, (LOAD_DATA_OUTER_LOOP_asn_10_itm[24:0]), {or_37_nl
      , and_196_nl , and_198_nl});
  assign mux_5_nl = MUX_s_1_2_2(or_1_cse, mux_4_cse, fsm_output[0]);
  assign dma_read_ctrl_write_reset_check_ResetChecker_dma_read_ctrl_write_reset_check_ResetChecker_and_nl
      = LOAD_DATA_INNER_LOOP_stage_0 & z_out_1_32;
  assign LOAD_DATA_OUTER_LOOP_mux_nl = MUX_s_1_2_2(dma_read_ctrl_write_reset_check_ResetChecker_dma_read_ctrl_write_reset_check_ResetChecker_and_nl,
      (~ z_out_1_32), and_dcpl_189);
  assign LOAD_DATA_OUTER_LOOP_mux_131_nl = MUX_v_32_2_2(offset_lpi_2, LOAD_BATCH_LOOP_b_sva,
      and_dcpl_214);
  assign not_116_nl = ~ and_dcpl_214;
  assign LOAD_DATA_OUTER_LOOP_LOAD_DATA_OUTER_LOOP_and_1_nl = MUX_v_25_2_2(25'b0000000000000000000000000,
      (LOAD_DATA_OUTER_LOOP_asn_10_itm[24:0]), not_116_nl);
  assign LOAD_DATA_OUTER_LOOP_mux_132_nl = MUX_v_7_2_2(LOAD_DATA_OUTER_LOOP_len_qr_6_0_lpi_2_dfm,
      7'b0000001, and_dcpl_214);
  assign nl_z_out = LOAD_DATA_OUTER_LOOP_mux_131_nl + ({LOAD_DATA_OUTER_LOOP_LOAD_DATA_OUTER_LOOP_and_1_nl
      , LOAD_DATA_OUTER_LOOP_mux_132_nl});
  assign z_out = nl_z_out[31:0];
  assign LOAD_BATCH_LOOP_mux1h_3_nl = MUX1HOT_v_32_6_2((~ (conf_info[63:32])), z_out,
      32'b00000000000000000000000010000001, ({16'b0000000000000000 , LOAD_DATA_INNER_LOOP_i_sva}),
      (~ (conf_info_crt_sva[31:0])), ({(~ z_out_2) , (~ (conf_info_crt_sva[6:0]))}),
      {and_dcpl_221 , and_dcpl_227 , and_dcpl_230 , and_dcpl_233 , and_dcpl_235 ,
      and_dcpl_238});
  assign LOAD_BATCH_LOOP_or_2_nl = (~(and_dcpl_221 | and_dcpl_230 | and_dcpl_235
      | and_dcpl_238)) | and_dcpl_227 | and_dcpl_233;
  assign LOAD_BATCH_LOOP_mux1h_4_nl = MUX1HOT_v_25_3_2((conf_info_crt_sva[63:39]),
      LOAD_DATA_OUTER_LOOP_s_31_7_sva, (LOAD_DATA_OUTER_LOOP_asn_10_itm[24:0]), {and_dcpl_227
      , and_dcpl_230 , and_dcpl_233});
  assign LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_nor_1_nl = ~(MUX_v_25_2_2(LOAD_BATCH_LOOP_mux1h_4_nl,
      25'b1111111111111111111111111, LOAD_BATCH_LOOP_or_1_ssc));
  assign LOAD_BATCH_LOOP_mux1h_5_nl = MUX1HOT_v_7_4_2(7'b0000001, (~ (conf_info_crt_sva[38:32])),
      (~ (conf_info_crt_sva[6:0])), (~ LOAD_DATA_OUTER_LOOP_len_qr_6_0_lpi_2_dfm),
      {LOAD_BATCH_LOOP_or_1_ssc , and_dcpl_227 , and_dcpl_230 , and_dcpl_233});
  assign nl_acc_1_nl = ({1'b1 , LOAD_BATCH_LOOP_mux1h_3_nl , LOAD_BATCH_LOOP_or_2_nl})
      + conv_u2u_33_34({LOAD_BATCH_LOOP_LOAD_BATCH_LOOP_nor_1_nl , LOAD_BATCH_LOOP_mux1h_5_nl
      , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[33:0];
  assign z_out_1_32 = readslicef_34_1_33(acc_1_nl);
  assign LOAD_DATA_INNER_LOOP_mux_127_nl = MUX_v_25_2_2(({9'b000000000 , LOAD_DATA_INNER_LOOP_i_sva}),
      LOAD_DATA_OUTER_LOOP_s_31_7_sva, and_dcpl_249);
  assign nl_z_out_2 = LOAD_DATA_INNER_LOOP_mux_127_nl + conv_s2u_2_25({and_dcpl_249
      , 1'b1});
  assign z_out_2 = nl_z_out_2[24:0];

  function automatic [24:0] MUX1HOT_v_25_3_2;
    input [24:0] input_2;
    input [24:0] input_1;
    input [24:0] input_0;
    input [2:0] sel;
    reg [24:0] result;
  begin
    result = input_0 & {25{sel[0]}};
    result = result | ( input_1 & {25{sel[1]}});
    result = result | ( input_2 & {25{sel[2]}});
    MUX1HOT_v_25_3_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_6_2;
    input [31:0] input_5;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [5:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    result = result | ( input_5 & {32{sel[5]}});
    MUX1HOT_v_32_6_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_126_2;
    input [6:0] input_125;
    input [6:0] input_124;
    input [6:0] input_123;
    input [6:0] input_122;
    input [6:0] input_121;
    input [6:0] input_120;
    input [6:0] input_119;
    input [6:0] input_118;
    input [6:0] input_117;
    input [6:0] input_116;
    input [6:0] input_115;
    input [6:0] input_114;
    input [6:0] input_113;
    input [6:0] input_112;
    input [6:0] input_111;
    input [6:0] input_110;
    input [6:0] input_109;
    input [6:0] input_108;
    input [6:0] input_107;
    input [6:0] input_106;
    input [6:0] input_105;
    input [6:0] input_104;
    input [6:0] input_103;
    input [6:0] input_102;
    input [6:0] input_101;
    input [6:0] input_100;
    input [6:0] input_99;
    input [6:0] input_98;
    input [6:0] input_97;
    input [6:0] input_96;
    input [6:0] input_95;
    input [6:0] input_94;
    input [6:0] input_93;
    input [6:0] input_92;
    input [6:0] input_91;
    input [6:0] input_90;
    input [6:0] input_89;
    input [6:0] input_88;
    input [6:0] input_87;
    input [6:0] input_86;
    input [6:0] input_85;
    input [6:0] input_84;
    input [6:0] input_83;
    input [6:0] input_82;
    input [6:0] input_81;
    input [6:0] input_80;
    input [6:0] input_79;
    input [6:0] input_78;
    input [6:0] input_77;
    input [6:0] input_76;
    input [6:0] input_75;
    input [6:0] input_74;
    input [6:0] input_73;
    input [6:0] input_72;
    input [6:0] input_71;
    input [6:0] input_70;
    input [6:0] input_69;
    input [6:0] input_68;
    input [6:0] input_67;
    input [6:0] input_66;
    input [6:0] input_65;
    input [6:0] input_64;
    input [6:0] input_63;
    input [6:0] input_62;
    input [6:0] input_61;
    input [6:0] input_60;
    input [6:0] input_59;
    input [6:0] input_58;
    input [6:0] input_57;
    input [6:0] input_56;
    input [6:0] input_55;
    input [6:0] input_54;
    input [6:0] input_53;
    input [6:0] input_52;
    input [6:0] input_51;
    input [6:0] input_50;
    input [6:0] input_49;
    input [6:0] input_48;
    input [6:0] input_47;
    input [6:0] input_46;
    input [6:0] input_45;
    input [6:0] input_44;
    input [6:0] input_43;
    input [6:0] input_42;
    input [6:0] input_41;
    input [6:0] input_40;
    input [6:0] input_39;
    input [6:0] input_38;
    input [6:0] input_37;
    input [6:0] input_36;
    input [6:0] input_35;
    input [6:0] input_34;
    input [6:0] input_33;
    input [6:0] input_32;
    input [6:0] input_31;
    input [6:0] input_30;
    input [6:0] input_29;
    input [6:0] input_28;
    input [6:0] input_27;
    input [6:0] input_26;
    input [6:0] input_25;
    input [6:0] input_24;
    input [6:0] input_23;
    input [6:0] input_22;
    input [6:0] input_21;
    input [6:0] input_20;
    input [6:0] input_19;
    input [6:0] input_18;
    input [6:0] input_17;
    input [6:0] input_16;
    input [6:0] input_15;
    input [6:0] input_14;
    input [6:0] input_13;
    input [6:0] input_12;
    input [6:0] input_11;
    input [6:0] input_10;
    input [6:0] input_9;
    input [6:0] input_8;
    input [6:0] input_7;
    input [6:0] input_6;
    input [6:0] input_5;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [125:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    result = result | ( input_3 & {7{sel[3]}});
    result = result | ( input_4 & {7{sel[4]}});
    result = result | ( input_5 & {7{sel[5]}});
    result = result | ( input_6 & {7{sel[6]}});
    result = result | ( input_7 & {7{sel[7]}});
    result = result | ( input_8 & {7{sel[8]}});
    result = result | ( input_9 & {7{sel[9]}});
    result = result | ( input_10 & {7{sel[10]}});
    result = result | ( input_11 & {7{sel[11]}});
    result = result | ( input_12 & {7{sel[12]}});
    result = result | ( input_13 & {7{sel[13]}});
    result = result | ( input_14 & {7{sel[14]}});
    result = result | ( input_15 & {7{sel[15]}});
    result = result | ( input_16 & {7{sel[16]}});
    result = result | ( input_17 & {7{sel[17]}});
    result = result | ( input_18 & {7{sel[18]}});
    result = result | ( input_19 & {7{sel[19]}});
    result = result | ( input_20 & {7{sel[20]}});
    result = result | ( input_21 & {7{sel[21]}});
    result = result | ( input_22 & {7{sel[22]}});
    result = result | ( input_23 & {7{sel[23]}});
    result = result | ( input_24 & {7{sel[24]}});
    result = result | ( input_25 & {7{sel[25]}});
    result = result | ( input_26 & {7{sel[26]}});
    result = result | ( input_27 & {7{sel[27]}});
    result = result | ( input_28 & {7{sel[28]}});
    result = result | ( input_29 & {7{sel[29]}});
    result = result | ( input_30 & {7{sel[30]}});
    result = result | ( input_31 & {7{sel[31]}});
    result = result | ( input_32 & {7{sel[32]}});
    result = result | ( input_33 & {7{sel[33]}});
    result = result | ( input_34 & {7{sel[34]}});
    result = result | ( input_35 & {7{sel[35]}});
    result = result | ( input_36 & {7{sel[36]}});
    result = result | ( input_37 & {7{sel[37]}});
    result = result | ( input_38 & {7{sel[38]}});
    result = result | ( input_39 & {7{sel[39]}});
    result = result | ( input_40 & {7{sel[40]}});
    result = result | ( input_41 & {7{sel[41]}});
    result = result | ( input_42 & {7{sel[42]}});
    result = result | ( input_43 & {7{sel[43]}});
    result = result | ( input_44 & {7{sel[44]}});
    result = result | ( input_45 & {7{sel[45]}});
    result = result | ( input_46 & {7{sel[46]}});
    result = result | ( input_47 & {7{sel[47]}});
    result = result | ( input_48 & {7{sel[48]}});
    result = result | ( input_49 & {7{sel[49]}});
    result = result | ( input_50 & {7{sel[50]}});
    result = result | ( input_51 & {7{sel[51]}});
    result = result | ( input_52 & {7{sel[52]}});
    result = result | ( input_53 & {7{sel[53]}});
    result = result | ( input_54 & {7{sel[54]}});
    result = result | ( input_55 & {7{sel[55]}});
    result = result | ( input_56 & {7{sel[56]}});
    result = result | ( input_57 & {7{sel[57]}});
    result = result | ( input_58 & {7{sel[58]}});
    result = result | ( input_59 & {7{sel[59]}});
    result = result | ( input_60 & {7{sel[60]}});
    result = result | ( input_61 & {7{sel[61]}});
    result = result | ( input_62 & {7{sel[62]}});
    result = result | ( input_63 & {7{sel[63]}});
    result = result | ( input_64 & {7{sel[64]}});
    result = result | ( input_65 & {7{sel[65]}});
    result = result | ( input_66 & {7{sel[66]}});
    result = result | ( input_67 & {7{sel[67]}});
    result = result | ( input_68 & {7{sel[68]}});
    result = result | ( input_69 & {7{sel[69]}});
    result = result | ( input_70 & {7{sel[70]}});
    result = result | ( input_71 & {7{sel[71]}});
    result = result | ( input_72 & {7{sel[72]}});
    result = result | ( input_73 & {7{sel[73]}});
    result = result | ( input_74 & {7{sel[74]}});
    result = result | ( input_75 & {7{sel[75]}});
    result = result | ( input_76 & {7{sel[76]}});
    result = result | ( input_77 & {7{sel[77]}});
    result = result | ( input_78 & {7{sel[78]}});
    result = result | ( input_79 & {7{sel[79]}});
    result = result | ( input_80 & {7{sel[80]}});
    result = result | ( input_81 & {7{sel[81]}});
    result = result | ( input_82 & {7{sel[82]}});
    result = result | ( input_83 & {7{sel[83]}});
    result = result | ( input_84 & {7{sel[84]}});
    result = result | ( input_85 & {7{sel[85]}});
    result = result | ( input_86 & {7{sel[86]}});
    result = result | ( input_87 & {7{sel[87]}});
    result = result | ( input_88 & {7{sel[88]}});
    result = result | ( input_89 & {7{sel[89]}});
    result = result | ( input_90 & {7{sel[90]}});
    result = result | ( input_91 & {7{sel[91]}});
    result = result | ( input_92 & {7{sel[92]}});
    result = result | ( input_93 & {7{sel[93]}});
    result = result | ( input_94 & {7{sel[94]}});
    result = result | ( input_95 & {7{sel[95]}});
    result = result | ( input_96 & {7{sel[96]}});
    result = result | ( input_97 & {7{sel[97]}});
    result = result | ( input_98 & {7{sel[98]}});
    result = result | ( input_99 & {7{sel[99]}});
    result = result | ( input_100 & {7{sel[100]}});
    result = result | ( input_101 & {7{sel[101]}});
    result = result | ( input_102 & {7{sel[102]}});
    result = result | ( input_103 & {7{sel[103]}});
    result = result | ( input_104 & {7{sel[104]}});
    result = result | ( input_105 & {7{sel[105]}});
    result = result | ( input_106 & {7{sel[106]}});
    result = result | ( input_107 & {7{sel[107]}});
    result = result | ( input_108 & {7{sel[108]}});
    result = result | ( input_109 & {7{sel[109]}});
    result = result | ( input_110 & {7{sel[110]}});
    result = result | ( input_111 & {7{sel[111]}});
    result = result | ( input_112 & {7{sel[112]}});
    result = result | ( input_113 & {7{sel[113]}});
    result = result | ( input_114 & {7{sel[114]}});
    result = result | ( input_115 & {7{sel[115]}});
    result = result | ( input_116 & {7{sel[116]}});
    result = result | ( input_117 & {7{sel[117]}});
    result = result | ( input_118 & {7{sel[118]}});
    result = result | ( input_119 & {7{sel[119]}});
    result = result | ( input_120 & {7{sel[120]}});
    result = result | ( input_121 & {7{sel[121]}});
    result = result | ( input_122 & {7{sel[122]}});
    result = result | ( input_123 & {7{sel[123]}});
    result = result | ( input_124 & {7{sel[124]}});
    result = result | ( input_125 & {7{sel[125]}});
    MUX1HOT_v_7_126_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_4_2;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [3:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    result = result | ( input_3 & {7{sel[3]}});
    MUX1HOT_v_7_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [24:0] MUX_v_25_2_2;
    input [24:0] input_0;
    input [24:0] input_1;
    input [0:0] sel;
    reg [24:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_25_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_34_1_33;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 33;
    readslicef_34_1_33 = tmp[0:0];
  end
  endfunction


  function automatic [24:0] conv_s2u_2_25 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_25 = {{23{vector[1]}}, vector};
  end
  endfunction


  function automatic [33:0] conv_u2u_33_34 ;
    input [32:0]  vector ;
  begin
    conv_u2u_33_34 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_store_output
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_store_output (
  clk, rst, conf_info, acc_done, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg,
      dma_write_chnl_val, dma_write_chnl_rdy, dma_write_chnl_msg, done, output_ready_channel_val,
      output_ready_channel_rdy, output_ready_channel_msg, plm_out_cns_dat, plm_out_cns_vld,
      plm_out_cns_rdy
);
  input clk;
  input rst;
  input [63:0] conf_info;
  output acc_done;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;
  input done;
  output output_ready_channel_val;
  input output_ready_channel_rdy;
  output output_ready_channel_msg;
  input [4095:0] plm_out_cns_dat;
  input plm_out_cns_vld;
  output plm_out_cns_rdy;


  // Interconnect Declarations
  wire STORE_MAIN_LOOP_plm_local_data_rsci_clken_d;
  wire [31:0] STORE_MAIN_LOOP_plm_local_data_rsci_d_d;
  wire [31:0] STORE_MAIN_LOOP_plm_local_data_rsci_q_d;
  wire [6:0] STORE_MAIN_LOOP_plm_local_data_rsci_radr_d;
  wire [6:0] STORE_MAIN_LOOP_plm_local_data_rsci_wadr_d;
  wire STORE_MAIN_LOOP_plm_local_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire STORE_MAIN_LOOP_plm_local_data_rsc_clken;
  wire [31:0] STORE_MAIN_LOOP_plm_local_data_rsc_q;
  wire [6:0] STORE_MAIN_LOOP_plm_local_data_rsc_radr;
  wire STORE_MAIN_LOOP_plm_local_data_rsc_we;
  wire [31:0] STORE_MAIN_LOOP_plm_local_data_rsc_d;
  wire [6:0] STORE_MAIN_LOOP_plm_local_data_rsc_wadr;
  wire STORE_MAIN_LOOP_plm_local_data_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  BLOCK_1R1W_RBW #(.addr_width(32'sd7),
  .data_width(32'sd32),
  .depth(32'sd128),
  .latency(32'sd1)) STORE_MAIN_LOOP_plm_local_data_rsc_comp (
      .clk(clk),
      .clken(STORE_MAIN_LOOP_plm_local_data_rsc_clken),
      .d(STORE_MAIN_LOOP_plm_local_data_rsc_d),
      .q(STORE_MAIN_LOOP_plm_local_data_rsc_q),
      .radr(STORE_MAIN_LOOP_plm_local_data_rsc_radr),
      .wadr(STORE_MAIN_LOOP_plm_local_data_rsc_wadr),
      .we(STORE_MAIN_LOOP_plm_local_data_rsc_we)
    );
  esp_acc_softmax_softmax_store_output_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_20_7_32_128_128_32_1_gen
      STORE_MAIN_LOOP_plm_local_data_rsci (
      .clken(STORE_MAIN_LOOP_plm_local_data_rsc_clken),
      .q(STORE_MAIN_LOOP_plm_local_data_rsc_q),
      .radr(STORE_MAIN_LOOP_plm_local_data_rsc_radr),
      .we(STORE_MAIN_LOOP_plm_local_data_rsc_we),
      .d(STORE_MAIN_LOOP_plm_local_data_rsc_d),
      .wadr(STORE_MAIN_LOOP_plm_local_data_rsc_wadr),
      .clken_d(STORE_MAIN_LOOP_plm_local_data_rsci_clken_d),
      .d_d(STORE_MAIN_LOOP_plm_local_data_rsci_d_d),
      .q_d(STORE_MAIN_LOOP_plm_local_data_rsci_q_d),
      .radr_d(STORE_MAIN_LOOP_plm_local_data_rsci_radr_d),
      .wadr_d(STORE_MAIN_LOOP_plm_local_data_rsci_wadr_d),
      .we_d(STORE_MAIN_LOOP_plm_local_data_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(STORE_MAIN_LOOP_plm_local_data_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(STORE_MAIN_LOOP_plm_local_data_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_softmax_softmax_store_output_store_output softmax_store_output_store_output_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .acc_done(acc_done),
      .dma_write_ctrl_val(dma_write_ctrl_val),
      .dma_write_ctrl_rdy(dma_write_ctrl_rdy),
      .dma_write_ctrl_msg(dma_write_ctrl_msg),
      .dma_write_chnl_val(dma_write_chnl_val),
      .dma_write_chnl_rdy(dma_write_chnl_rdy),
      .dma_write_chnl_msg(dma_write_chnl_msg),
      .done(done),
      .output_ready_channel_val(output_ready_channel_val),
      .output_ready_channel_rdy(output_ready_channel_rdy),
      .output_ready_channel_msg(output_ready_channel_msg),
      .plm_out_cns_dat(plm_out_cns_dat),
      .plm_out_cns_vld(plm_out_cns_vld),
      .plm_out_cns_rdy(plm_out_cns_rdy),
      .STORE_MAIN_LOOP_plm_local_data_rsci_clken_d(STORE_MAIN_LOOP_plm_local_data_rsci_clken_d),
      .STORE_MAIN_LOOP_plm_local_data_rsci_d_d(STORE_MAIN_LOOP_plm_local_data_rsci_d_d),
      .STORE_MAIN_LOOP_plm_local_data_rsci_q_d(STORE_MAIN_LOOP_plm_local_data_rsci_q_d),
      .STORE_MAIN_LOOP_plm_local_data_rsci_radr_d(STORE_MAIN_LOOP_plm_local_data_rsci_radr_d),
      .STORE_MAIN_LOOP_plm_local_data_rsci_wadr_d(STORE_MAIN_LOOP_plm_local_data_rsci_wadr_d),
      .STORE_MAIN_LOOP_plm_local_data_rsci_readA_r_ram_ir_internal_RMASK_B_d(STORE_MAIN_LOOP_plm_local_data_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .STORE_MAIN_LOOP_plm_local_data_rsci_we_d_pff(STORE_MAIN_LOOP_plm_local_data_rsci_we_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_compute_kernel
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_compute_kernel (
  clk, rst, conf_info, done, input_ready_channel_val, input_ready_channel_rdy, input_ready_channel_msg,
      output_ready_channel_val, output_ready_channel_rdy, output_ready_channel_msg,
      plm_in_cns_dat, plm_in_cns_vld, plm_in_cns_rdy, plm_out_cns_dat, plm_out_cns_vld,
      plm_out_cns_rdy
);
  input clk;
  input rst;
  input [63:0] conf_info;
  input done;
  output input_ready_channel_val;
  input input_ready_channel_rdy;
  output input_ready_channel_msg;
  input output_ready_channel_val;
  output output_ready_channel_rdy;
  input output_ready_channel_msg;
  input [4095:0] plm_in_cns_dat;
  input plm_in_cns_vld;
  output plm_in_cns_rdy;
  output [4095:0] plm_out_cns_dat;
  output plm_out_cns_vld;
  input plm_out_cns_rdy;


  // Interconnect Declarations
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_adra_d;
  wire [2047:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_da_d;
  wire [2047:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_wea_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_adra_d;
  wire [2047:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_da_d;
  wire [2047:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_wea_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_adra_d;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_da_d;
  wire [2047:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_wea_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_adra_d;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_da_d;
  wire [2047:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_wea_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [1:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  wire [93:0] CALC_SOFTMAX_LOOP_mul_cmp_b;
  wire [94:0] CALC_SOFTMAX_LOOP_mul_cmp_z;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_clken;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_q;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_radr;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_we;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_d;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wadr;
  wire COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_clkb_en;
  wire COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_clka_en;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_qb;
  wire COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_web;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_db;
  wire COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_adrb;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_qa;
  wire COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_wea;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_da;
  wire COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_adra;
  wire COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_clkb_en;
  wire COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_clka_en;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_qb;
  wire COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_web;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_db;
  wire COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_adrb;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_qa;
  wire COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_wea;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_da;
  wire COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_adra;
  wire COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_clkb_en;
  wire COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_clka_en;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_qb;
  wire COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_web;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_db;
  wire COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_adrb;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_qa;
  wire COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_wea;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_da;
  wire COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_adra;
  wire COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_clkb_en;
  wire COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_clka_en;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_qb;
  wire COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_web;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_db;
  wire COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_adrb;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_qa;
  wire COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_wea;
  wire [1023:0] COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_da;
  wire COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_adra;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [2047:0] nl_COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_da_d;
  assign nl_COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_da_d = {COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_da_d
      , {512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
      , 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000}};
  wire [2047:0] nl_COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_da_d;
  assign nl_COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_da_d = {COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_da_d
      , {512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
      , 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000}};
  esp_acc_softmax_mgc_mul_pipe #(.width_a(32'sd67),
  .signd_a(32'sd0),
  .width_b(32'sd94),
  .signd_b(32'sd0),
  .width_z(32'sd95),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) CALC_SOFTMAX_LOOP_mul_cmp (
      .a(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d),
      .b(CALC_SOFTMAX_LOOP_mul_cmp_b),
      .clk(clk),
      .en(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(CALC_SOFTMAX_LOOP_mul_cmp_z)
    );
  BLOCK_1R1W_RBW #(.addr_width(32'sd7),
  .data_width(32'sd67),
  .depth(32'sd128),
  .latency(32'sd1)) ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_comp
      (
      .clk(clk),
      .clken(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_clken),
      .d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_d),
      .q(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_q),
      .radr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_radr),
      .wadr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wadr),
      .we(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_we)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd1),
  .data_width(32'sd1024),
  .depth(32'sd2),
  .latency(32'sd1)) COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_comp (
      .adra(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_adra),
      .adrb(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_adrb),
      .clka(clk),
      .clka_en(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_clkb_en),
      .clkb(clk),
      .clkb_en(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_clkb_en),
      .da(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_da),
      .db(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_db),
      .qa(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_qa),
      .qb(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_qb),
      .wea(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_wea),
      .web(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd1),
  .data_width(32'sd1024),
  .depth(32'sd2),
  .latency(32'sd1)) COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_comp (
      .adra(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_adra),
      .adrb(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_adrb),
      .clka(clk),
      .clka_en(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_clkb_en),
      .clkb(clk),
      .clkb_en(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_clkb_en),
      .da(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_da),
      .db(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_db),
      .qa(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_qa),
      .qb(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_qb),
      .wea(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_wea),
      .web(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd1),
  .data_width(32'sd1024),
  .depth(32'sd2),
  .latency(32'sd1)) COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_comp (
      .adra(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_adra),
      .adrb(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_adrb),
      .clka(clk),
      .clka_en(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_clkb_en),
      .clkb(clk),
      .clkb_en(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_clkb_en),
      .da(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_da),
      .db(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_db),
      .qa(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_qa),
      .qb(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_qb),
      .wea(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_wea),
      .web(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd1),
  .data_width(32'sd1024),
  .depth(32'sd2),
  .latency(32'sd1)) COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_comp (
      .adra(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_adra),
      .adrb(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_adrb),
      .clka(clk),
      .clka_en(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_clkb_en),
      .clkb(clk),
      .clkb_en(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_clkb_en),
      .da(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_da),
      .db(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_db),
      .qa(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_qa),
      .qb(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_qb),
      .wea(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_wea),
      .web(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_web)
    );
  esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_19_7_67_128_128_67_1_gen
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci
      (
      .clken(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_clken),
      .q(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_q),
      .radr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_radr),
      .we(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_we),
      .d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_d),
      .wadr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wadr),
      .clken_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d),
      .d_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d),
      .q_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d),
      .radr_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d),
      .wadr_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d),
      .we_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_48_1_1024_2_2_1024_1_gen
      COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i (
      .clkb_en(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_clkb_en),
      .clka_en(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_clka_en),
      .qb(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_qb),
      .web(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_web),
      .db(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_db),
      .adrb(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_adrb),
      .qa(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_qa),
      .wea(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_wea),
      .da(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_da),
      .adra(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_adra),
      .adra_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_adra_d),
      .clka(clk),
      .clka_en_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d),
      .clkb_en_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d),
      .da_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_da_d),
      .qa_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d),
      .wea_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_wea_d),
      .rwA_rw_ram_ir_internal_RMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d)
    );
  esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_49_1_1024_2_2_1024_1_gen
      COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i (
      .clkb_en(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_clkb_en),
      .clka_en(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_clka_en),
      .qb(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_qb),
      .web(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_web),
      .db(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_db),
      .adrb(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_adrb),
      .qa(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_qa),
      .wea(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_wea),
      .da(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_da),
      .adra(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_adra),
      .adra_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_adra_d),
      .clka(clk),
      .clka_en_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d),
      .clkb_en_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d),
      .da_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_da_d),
      .qa_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d),
      .wea_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_wea_d),
      .rwA_rw_ram_ir_internal_RMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d)
    );
  esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_50_1_1024_2_2_1024_1_gen
      COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i (
      .clkb_en(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_clkb_en),
      .clka_en(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_clka_en),
      .qb(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_qb),
      .web(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_web),
      .db(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_db),
      .adrb(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_adrb),
      .qa(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_qa),
      .wea(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_wea),
      .da(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_da),
      .adra(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_adra),
      .adra_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_adra_d),
      .clka(clk),
      .clka_en_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d),
      .clkb_en_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d),
      .da_d(nl_COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_da_d[2047:0]),
      .qa_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d),
      .wea_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_wea_d),
      .rwA_rw_ram_ir_internal_RMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d)
    );
  esp_acc_softmax_softmax_compute_kernel_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_51_1_1024_2_2_1024_1_gen
      COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i (
      .clkb_en(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_clkb_en),
      .clka_en(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_clka_en),
      .qb(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_qb),
      .web(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_web),
      .db(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_db),
      .adrb(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_adrb),
      .qa(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_qa),
      .wea(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_wea),
      .da(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_da),
      .adra(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_adra),
      .adra_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_adra_d),
      .clka(clk),
      .clka_en_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d),
      .clkb_en_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d),
      .da_d(nl_COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_da_d[2047:0]),
      .qa_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d),
      .wea_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_wea_d),
      .rwA_rw_ram_ir_internal_RMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d)
    );
  esp_acc_softmax_softmax_compute_kernel_compute_kernel softmax_compute_kernel_compute_kernel_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .done(done),
      .input_ready_channel_val(input_ready_channel_val),
      .input_ready_channel_rdy(input_ready_channel_rdy),
      .input_ready_channel_msg(input_ready_channel_msg),
      .output_ready_channel_val(output_ready_channel_val),
      .output_ready_channel_rdy(output_ready_channel_rdy),
      .output_ready_channel_msg(output_ready_channel_msg),
      .plm_in_cns_dat(plm_in_cns_dat),
      .plm_in_cns_vld(plm_in_cns_vld),
      .plm_in_cns_rdy(plm_in_cns_rdy),
      .plm_out_cns_dat(plm_out_cns_dat),
      .plm_out_cns_vld(plm_out_cns_vld),
      .plm_out_cns_rdy(plm_out_cns_rdy),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_clken_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_adra_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_adra_d),
      .COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_da_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_da_d),
      .COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_qa_d),
      .COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_wea_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_wea_d),
      .COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d),
      .COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_adra_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_adra_d),
      .COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_da_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_da_d),
      .COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_qa_d),
      .COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_wea_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_wea_d),
      .COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_in_data_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d),
      .COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_adra_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_adra_d),
      .COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_da_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_da_d),
      .COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_qa_d),
      .COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_wea_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_wea_d),
      .COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d),
      .COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_adra_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_adra_d),
      .COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_da_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_da_d),
      .COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_qa_d),
      .COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_wea_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_wea_d),
      .COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d(COMPUTE_OUTER_LOOP_plm_local_out_data_rsc_0_1_i_rwA_rw_ram_ir_internal_WMASK_B_d),
      .CALC_SOFTMAX_LOOP_mul_cmp_b(CALC_SOFTMAX_LOOP_mul_cmp_b),
      .CALC_SOFTMAX_LOOP_mul_cmp_z(CALC_SOFTMAX_LOOP_mul_cmp_z),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_softmax_load_input
// ------------------------------------------------------------------


module esp_acc_softmax_softmax_load_input (
  clk, rst, conf_info, dma_read_ctrl_val, dma_read_ctrl_rdy, dma_read_ctrl_msg, dma_read_chnl_val,
      dma_read_chnl_rdy, dma_read_chnl_msg, done, input_ready_channel_val, input_ready_channel_rdy,
      input_ready_channel_msg, plm_in_cns_dat, plm_in_cns_vld, plm_in_cns_rdy
);
  input clk;
  input rst;
  input [63:0] conf_info;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  input done;
  input input_ready_channel_val;
  output input_ready_channel_rdy;
  input input_ready_channel_msg;
  output [4095:0] plm_in_cns_dat;
  output plm_in_cns_vld;
  input plm_in_cns_rdy;


  // Interconnect Declarations
  wire LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_clken_d;
  wire [31:0] LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_d_d;
  wire [31:0] LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d;
  wire [6:0] LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_radr_d;
  wire [6:0] LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_wadr_d;
  wire LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_clken;
  wire [31:0] LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_q;
  wire [6:0] LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_radr;
  wire LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_we;
  wire [31:0] LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_d;
  wire [6:0] LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_wadr;
  wire LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  BLOCK_1R1W_RBW #(.addr_width(32'sd7),
  .data_width(32'sd32),
  .depth(32'sd128),
  .latency(32'sd1)) LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_comp (
      .clk(clk),
      .clken(LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_clken),
      .d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_d),
      .q(LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_q),
      .radr(LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_radr),
      .wadr(LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_wadr),
      .we(LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_we)
    );
  esp_acc_softmax_softmax_load_input_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_16_7_32_128_128_32_1_gen
      LOAD_DATA_OUTER_LOOP_plm_local_data_rsci (
      .clken(LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_clken),
      .q(LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_q),
      .radr(LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_radr),
      .we(LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_we),
      .d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_d),
      .wadr(LOAD_DATA_OUTER_LOOP_plm_local_data_rsc_wadr),
      .clken_d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_clken_d),
      .d_d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_d_d),
      .q_d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d),
      .radr_d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_radr_d),
      .wadr_d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_wadr_d),
      .we_d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_softmax_softmax_load_input_load_input softmax_load_input_load_input_inst
      (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .dma_read_ctrl_val(dma_read_ctrl_val),
      .dma_read_ctrl_rdy(dma_read_ctrl_rdy),
      .dma_read_ctrl_msg(dma_read_ctrl_msg),
      .dma_read_chnl_val(dma_read_chnl_val),
      .dma_read_chnl_rdy(dma_read_chnl_rdy),
      .dma_read_chnl_msg(dma_read_chnl_msg),
      .done(done),
      .input_ready_channel_val(input_ready_channel_val),
      .input_ready_channel_rdy(input_ready_channel_rdy),
      .input_ready_channel_msg(input_ready_channel_msg),
      .plm_in_cns_dat(plm_in_cns_dat),
      .plm_in_cns_vld(plm_in_cns_vld),
      .plm_in_cns_rdy(plm_in_cns_rdy),
      .LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_clken_d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_clken_d),
      .LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_d_d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_d_d),
      .LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_q_d),
      .LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_radr_d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_radr_d),
      .LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_wadr_d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_wadr_d),
      .LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_readA_r_ram_ir_internal_RMASK_B_d(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_we_d_pff(LOAD_DATA_OUTER_LOOP_plm_local_data_rsci_we_d_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    softmax_basic_fx32_dma64
// ------------------------------------------------------------------


module softmax_basic_fx32_dma64 (
  clk, rst, conf_info, conf_done, acc_done, debug, dma_read_ctrl_val, dma_read_ctrl_rdy,
      dma_read_ctrl_msg, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg,
      dma_read_chnl_val, dma_read_chnl_rdy, dma_read_chnl_msg, dma_write_chnl_val,
      dma_write_chnl_rdy, dma_write_chnl_msg
);
  input clk;
  input rst;
  input [63:0] conf_info;
  input conf_done;
  output acc_done;
  output [31:0] debug;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;


  // Interconnect Declarations
  wire done;
  wire input_ready_channel_val;
  wire input_ready_channel_rdy;
  wire input_ready_channel_msg;
  wire output_ready_channel_val;
  wire output_ready_channel_rdy;
  wire output_ready_channel_msg;
  wire [4095:0] plm_in_cns_dat_nsoftmax_load_input_inst;
  wire plm_in_cns_rdy_nsoftmax_load_input_inst;
  wire [4095:0] plm_in_cns_dat_nsoftmax_compute_kernel_inst;
  wire plm_in_cns_vld_nsoftmax_compute_kernel_inst;
  wire [4095:0] plm_out_cns_dat_nsoftmax_compute_kernel_inst;
  wire plm_out_cns_rdy_nsoftmax_compute_kernel_inst;
  wire [4095:0] plm_out_cns_dat_nsoftmax_store_output_inst;
  wire plm_out_cns_vld_nsoftmax_store_output_inst;
  wire plm_in_cns_vld_nsoftmax_load_input_inst_bud;
  wire plm_in_cns_rdy_nsoftmax_compute_kernel_inst_bud;
  wire plm_out_cns_vld_nsoftmax_compute_kernel_inst_bud;
  wire plm_out_cns_rdy_nsoftmax_store_output_inst_bud;
  wire plm_in_unc_2;
  wire plm_in_idle;
  wire plm_out_unc_2;
  wire plm_out_idle;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_ccs_pipe_v5 #(.rscid(32'sd25),
  .width(32'sd4096),
  .sz_width(32'sd1),
  .fifo_sz(32'sd32),
  .log2_sz(32'sd5),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) plm_in_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(1'b1),
      .srst(rst),
      .din_rdy(plm_in_cns_rdy_nsoftmax_load_input_inst),
      .din_vld(plm_in_cns_vld_nsoftmax_load_input_inst_bud),
      .din(plm_in_cns_dat_nsoftmax_load_input_inst),
      .dout_rdy(plm_in_cns_rdy_nsoftmax_compute_kernel_inst_bud),
      .dout_vld(plm_in_cns_vld_nsoftmax_compute_kernel_inst),
      .dout(plm_in_cns_dat_nsoftmax_compute_kernel_inst),
      .sz(plm_in_unc_2),
      .sz_req(1'b0),
      .is_idle(plm_in_idle)
    );
  esp_acc_softmax_ccs_pipe_v5 #(.rscid(32'sd26),
  .width(32'sd4096),
  .sz_width(32'sd1),
  .fifo_sz(32'sd32),
  .log2_sz(32'sd5),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) plm_out_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(1'b1),
      .srst(rst),
      .din_rdy(plm_out_cns_rdy_nsoftmax_compute_kernel_inst),
      .din_vld(plm_out_cns_vld_nsoftmax_compute_kernel_inst_bud),
      .din(plm_out_cns_dat_nsoftmax_compute_kernel_inst),
      .dout_rdy(plm_out_cns_rdy_nsoftmax_store_output_inst_bud),
      .dout_vld(plm_out_cns_vld_nsoftmax_store_output_inst),
      .dout(plm_out_cns_dat_nsoftmax_store_output_inst),
      .sz(plm_out_unc_2),
      .sz_req(1'b0),
      .is_idle(plm_out_idle)
    );
  esp_acc_softmax_softmax_load_input softmax_load_input_inst (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .dma_read_ctrl_val(dma_read_ctrl_val),
      .dma_read_ctrl_rdy(dma_read_ctrl_rdy),
      .dma_read_ctrl_msg(dma_read_ctrl_msg),
      .dma_read_chnl_val(dma_read_chnl_val),
      .dma_read_chnl_rdy(dma_read_chnl_rdy),
      .dma_read_chnl_msg(dma_read_chnl_msg),
      .done(done),
      .input_ready_channel_val(input_ready_channel_val),
      .input_ready_channel_rdy(input_ready_channel_rdy),
      .input_ready_channel_msg(input_ready_channel_msg),
      .plm_in_cns_dat(plm_in_cns_dat_nsoftmax_load_input_inst),
      .plm_in_cns_vld(plm_in_cns_vld_nsoftmax_load_input_inst_bud),
      .plm_in_cns_rdy(plm_in_cns_rdy_nsoftmax_load_input_inst)
    );
  esp_acc_softmax_softmax_compute_kernel softmax_compute_kernel_inst (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .done(done),
      .input_ready_channel_val(input_ready_channel_val),
      .input_ready_channel_rdy(input_ready_channel_rdy),
      .input_ready_channel_msg(input_ready_channel_msg),
      .output_ready_channel_val(output_ready_channel_val),
      .output_ready_channel_rdy(output_ready_channel_rdy),
      .output_ready_channel_msg(output_ready_channel_msg),
      .plm_in_cns_dat(plm_in_cns_dat_nsoftmax_compute_kernel_inst),
      .plm_in_cns_vld(plm_in_cns_vld_nsoftmax_compute_kernel_inst),
      .plm_in_cns_rdy(plm_in_cns_rdy_nsoftmax_compute_kernel_inst_bud),
      .plm_out_cns_dat(plm_out_cns_dat_nsoftmax_compute_kernel_inst),
      .plm_out_cns_vld(plm_out_cns_vld_nsoftmax_compute_kernel_inst_bud),
      .plm_out_cns_rdy(plm_out_cns_rdy_nsoftmax_compute_kernel_inst)
    );
  esp_acc_softmax_softmax_store_output softmax_store_output_inst (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .acc_done(acc_done),
      .dma_write_ctrl_val(dma_write_ctrl_val),
      .dma_write_ctrl_rdy(dma_write_ctrl_rdy),
      .dma_write_ctrl_msg(dma_write_ctrl_msg),
      .dma_write_chnl_val(dma_write_chnl_val),
      .dma_write_chnl_rdy(dma_write_chnl_rdy),
      .dma_write_chnl_msg(dma_write_chnl_msg),
      .done(done),
      .output_ready_channel_val(output_ready_channel_val),
      .output_ready_channel_rdy(output_ready_channel_rdy),
      .output_ready_channel_msg(output_ready_channel_msg),
      .plm_out_cns_dat(plm_out_cns_dat_nsoftmax_store_output_inst),
      .plm_out_cns_vld(plm_out_cns_vld_nsoftmax_store_output_inst),
      .plm_out_cns_rdy(plm_out_cns_rdy_nsoftmax_store_output_inst_bud)
    );
  esp_acc_softmax_softmax_config_accelerator softmax_config_accelerator_inst (
      .clk(clk),
      .rst(rst),
      .conf_done(conf_done),
      .done(done)
    );
endmodule



