
//------> ./softmax_sysc_Connections_OutBlockingless_dma_info_tcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_sysc_Connections_OutBlockingless_dma_info_tcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_sysc_Connections_OutBlockingless_dma_info_tcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue Jun  9 14:16:35 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core
    (
  this_val, this_rdy, this_msg, m_index_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [66:0] this_msg;
  input [31:0] m_index_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire [31:0] m_index_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [24:0] m_index_slc_m_index_31_7_psp_lpi_1_dfm;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  reg reg_C_35_1_reg_32;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd32)) m_index_rsci (
      .dat(m_index_rsc_dat),
      .idat(m_index_rsci_idat)
    );
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 #(.rscid(32'sd19),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 #(.rscid(32'sd22)) ccs_ccore_done_synci
      (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign this_msg = {1'b0 , ({{1{reg_C_35_1_reg_32}}, reg_C_35_1_reg_32}) , 24'b000000000000000000000000
      , reg_C_35_1_reg_32 , 7'b0000000 , m_index_slc_m_index_31_7_psp_lpi_1_dfm ,
      7'b0000000};
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_val <= 1'b0;
    end
    else if ( or_4_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      reg_C_35_1_reg_32 <= 1'b0;
    end
    else if ( (~((~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1) | this_rdy)) | ccs_ccore_start_rsci_idat
        ) begin
      reg_C_35_1_reg_32 <= 1'b1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      m_index_slc_m_index_31_7_psp_lpi_1_dfm <= 25'b0000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      m_index_slc_m_index_31_7_psp_lpi_1_dfm <= m_index_rsci_idat[31:7];
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_index_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  input this_rdy;
  output [66:0] this_msg;
  input [31:0] m_index_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push_core_inst (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_index_rsc_dat(m_index_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_sysc_Connections_InBlockingless_dma_data_tcomma_Connections_SYN_PORTgreater_Pop_mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ./softmax_sysc_Connections_InBlockingless_dma_data_tcomma_Connections_SYN_PORTgreater_Pop_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_sysc_Connections_InBlockingless_dma_data_tcomma_Connections_SYN_PORTgreater_Pop_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_sysc_Connections_InBlockingless_dma_data_tcomma_Connections_SYN_PORTgreater_Pop.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue Jun  9 14:16:34 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_Connections_InBlocking_dma_data_t_Connections_SYN_PORT_Pop_core
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_Connections_InBlocking_dma_data_t_Connections_SYN_PORT_Pop_core
    (
  this_val, this_rdy, this_msg, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [63:0] this_msg;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_2_cse;
  wire this_rdy_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [63:0] nl_return_rsci_d;
  assign nl_return_rsci_d = this_msg;
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_val;
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_mgc_out_dreg_v2 #(.rscid(32'sd4),
  .width(32'sd64)) return_rsci (
      .d(nl_return_rsci_d[63:0]),
      .z(return_rsc_z)
    );
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 #(.rscid(32'sd18),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 #(.rscid(32'sd21)) ccs_ccore_done_synci
      (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign or_2_cse = ccs_ccore_start_rsci_idat | (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_val));
  assign this_rdy_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_val
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_rdy <= 1'b0;
    end
    else if ( or_2_cse | this_rdy_mx0c1 ) begin
      this_rdy <= ~ this_rdy_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_2_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_dma_data_t_Connections_SYN_PORT_Pop
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_Connections_InBlocking_dma_data_t_Connections_SYN_PORT_Pop (
  this_val, this_rdy, this_msg, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  input this_val;
  output this_rdy;
  input [63:0] this_msg;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_Connections_InBlocking_dma_data_t_Connections_SYN_PORT_Pop_core
      Connections_InBlocking_dma_data_t_Connections_SYN_PORT_Pop_core_inst (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_sysc_Connections_OutBlockingless_dma_data_tcomma_Connections_SYN_PORTgreater_Push_ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ./softmax_sysc_Connections_OutBlockingless_dma_data_tcomma_Connections_SYN_PORTgreater_Push_ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ./softmax_sysc_Connections_OutBlockingless_dma_data_tcomma_Connections_SYN_PORTgreater_Push.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue Jun  9 14:16:31 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_Connections_OutBlocking_dma_data_t_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_esp_acc_softmax_sysc_Connections_OutBlocking_dma_data_t_Connections_SYN_PORT_Push_core
    (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [63:0] this_msg;
  input [63:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;


  // Interconnect Declarations
  wire [63:0] m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg [31:0] m_slc_m_31_0_psp_lpi_1_dfm;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_4_cse;
  reg reg_C_32_11011110101011011011111011101111_1_reg_30;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd64)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_in_v1 #(.rscid(32'sd17),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_ccs_sync_out_vld_v1 #(.rscid(32'sd20)) ccs_ccore_done_synci
      (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign this_msg = signext_64_63({reg_C_32_11011110101011011011111011101111_1_reg_30
      , 1'b0 , ({{3{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , reg_C_32_11011110101011011011111011101111_1_reg_30 , 1'b0 , reg_C_32_11011110101011011011111011101111_1_reg_30
      , 1'b0 , ({{1{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{1{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{4{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{2{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , 1'b0 , ({{3{reg_C_32_11011110101011011011111011101111_1_reg_30}}, reg_C_32_11011110101011011011111011101111_1_reg_30})
      , m_slc_m_31_0_psp_lpi_1_dfm});
  assign or_4_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      this_val <= 1'b0;
    end
    else if ( or_4_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      reg_C_32_11011110101011011011111011101111_1_reg_30 <= 1'b0;
    end
    else if ( (~((~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1) | this_rdy)) | ccs_ccore_start_rsci_idat
        ) begin
      reg_C_32_11011110101011011011111011101111_1_reg_30 <= 1'b1;
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      m_slc_m_31_0_psp_lpi_1_dfm <= 32'b00000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      m_slc_m_31_0_psp_lpi_1_dfm <= m_rsci_idat[31:0];
    end
  end
  always @(posedge ccs_MIO_clk) begin
    if ( ~ ccs_MIO_srst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_4_cse;
    end
  end

  function automatic [63:0] signext_64_63;
    input [62:0] vector;
  begin
    signext_64_63= {{1{vector[62]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_dma_data_t_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_Connections_OutBlocking_dma_data_t_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_srst
);
  output this_val;
  input this_rdy;
  output [63:0] this_msg;
  input [63:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_srst;



  // Interconnect Declarations for Component Instantiations
  esp_acc_softmax_sysc_esp_acc_softmax_sysc_Connections_OutBlocking_dma_data_t_Connections_SYN_PORT_Push_core
      Connections_OutBlocking_dma_data_t_Connections_SYN_PORT_Push_core_inst (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_rsc_dat(m_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_srst(ccs_MIO_srst)
    );
endmodule




//------> ./softmax_sysc_mgc_mul_pipe_beh.v 
//
// File:      $Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v
//
// BASELINE:  Catapult-C version 2006b.63
// MODIFIED:  2007-04-03, tnagler
//
// Note: this file uses Verilog2001 features;
//       please enable Verilog2001 in the flow!

module esp_acc_softmax_sysc_mgc_mul_pipe (a, b, clk, en, a_rst, s_rst, z);

    // Parameters:
    parameter integer width_a = 32'd4;  // input a bit width
    parameter         signd_a =  1'b1;  // input a type (1=signed, 0=unsigned)
    parameter integer width_b = 32'd4;  // input b bit width
    parameter         signd_b =  1'b1;  // input b type (1=signed, 0=unsigned)
    parameter integer width_z = 32'd8;  // result bit width (= width_a + width_b)
    parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
    parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
    parameter    a_rst_active =  1'b1;  // unused
    parameter    s_rst_active =  1'b1;  // unused
    parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
    parameter integer n_inreg = 32'd0;  // number of input registers

    localparam integer width_ab = width_a + width_b;  // multiplier result width
    localparam integer n_inreg_min = (n_inreg > 1) ? (n_inreg-1) : 0; // for Synopsys DC

    // I/O ports:
    input  [width_a-1:0] a;      // input A
    input  [width_b-1:0] b;      // input B
    input                clk;    // clock
    input                en;     // enable
    input                a_rst;  // async reset (unused)
    input                s_rst;  // sync reset (unused)
    output [width_z-1:0] z;      // output


    // Input registers:

    wire [width_a-1:0] a_f;
    wire [width_b-1:0] b_f;

    integer i;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(negedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i];
                    b_reg[i+1] <= b_reg[i];
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    else
    begin: POS_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a,
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(posedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i];
                    b_reg[i+1] <= b_reg[i];
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    endgenerate


    // Output:
    wire [width_z-1:0]  xz;

    function signed [width_z-1:0] conv_signed;
      input signed [width_ab-1:0] res;
      conv_signed = res[width_z-1:0];
    endfunction

    generate
      wire signed [width_ab-1:0] res;
      if ( (signd_a == 1'b1) && (signd_b == 1'b1) )
      begin: SIGNED_AB
              assign res = $signed(a_f) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b1) && (signd_b == 1'b0) )
      begin: SIGNED_A
              assign res = $signed(a_f) * $signed({1'b0, b_f});
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b0) && (signd_b == 1'b1) )
      begin: SIGNED_B
              assign res = $signed({1'b0,a_f}) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else
      begin: UNSIGNED_AB
              assign res = a_f * b_f;
	      assign xz = res[width_z-1:0];
      end
    endgenerate


    // Output registers:

    reg  [width_z-1:0] reg_array[stages-2:0];
    wire [width_z-1:0] z;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE2
        always @(negedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz;
                else
                    reg_array[i] <= reg_array[i-1];
    end
    else
    begin: POS_EDGE2
        always @(posedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz;
                else
                    reg_array[i] <= reg_array[i-1];
    end
    endgenerate

    assign z = reg_array[stages-2];
endmodule

//------> ./softmax_sysc_mgc_shift_br_beh_v5.v 
module esp_acc_softmax_sysc_mgc_shift_br_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_s(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_s(a,s,1'b0);
     end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshr_u

   //Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction

endmodule

//------> ./softmax_sysc_mgc_shift_bl_beh_v5.v 
module esp_acc_softmax_sysc_mgc_shift_bl_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate if ( signd_a )
   begin: SGNED
     assign z = fshl_s(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
     assign z = fshl_s(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

endmodule

//------> ./softmax_sysc_mgc_shift_l_beh_v5.v 
module esp_acc_softmax_sysc_mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./softmax_sysc_leading_sign_74_0.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
//
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue Jun  9 14:16:33 2020
// ----------------------------------------------------------------------

//
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_74_0
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_leading_sign_74_0 (
  mantissa, rtn
);
  input [73:0] mantissa;
  output [6:0] rtn;


  // Interconnect Declarations
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_24;
  wire c_h_1_27;
  wire c_h_1_28;
  wire c_h_1_29;
  wire c_h_1_30;
  wire c_h_1_33;
  wire c_h_1_34;
  wire c_h_1_35;
  wire ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc;

  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_1_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_292_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_2_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_or_2_nl;
  wire[0:0] ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_nor_nl;

  // Interconnect Declarations for Component Instantiations
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2
      = ~((mantissa[71:70]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1
      = ~((mantissa[73:72]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1
      = ~((mantissa[69:68]!=2'b00));
  assign c_h_1_2 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3
      = (mantissa[67:66]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2
      = ~((mantissa[63:62]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1
      = ~((mantissa[65:64]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1
      = ~((mantissa[61:60]!=2'b00));
  assign c_h_1_5 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4
      = (mantissa[59:58]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1
      & c_h_1_5;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2
      = ~((mantissa[55:54]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1
      = ~((mantissa[57:56]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1
      = ~((mantissa[53:52]!=2'b00));
  assign c_h_1_9 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3
      = (mantissa[51:50]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2
      = ~((mantissa[47:46]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1
      = ~((mantissa[49:48]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1
      = ~((mantissa[45:44]!=2'b00));
  assign c_h_1_12 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5
      = (mantissa[43:42]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1
      & c_h_1_12 & c_h_1_13;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2
      = ~((mantissa[39:38]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1
      = ~((mantissa[41:40]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1
      = ~((mantissa[37:36]!=2'b00));
  assign c_h_1_17 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3
      = (mantissa[35:34]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2
      = ~((mantissa[31:30]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1
      = ~((mantissa[33:32]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1
      = ~((mantissa[29:28]!=2'b00));
  assign c_h_1_20 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4
      = (mantissa[27:26]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1
      & c_h_1_20;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2
      = ~((mantissa[23:22]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1
      = ~((mantissa[25:24]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1
      = ~((mantissa[21:20]!=2'b00));
  assign c_h_1_24 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3
      = (mantissa[19:18]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2
      = ~((mantissa[15:14]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1
      = ~((mantissa[17:16]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1
      = ~((mantissa[13:12]!=2'b00));
  assign c_h_1_27 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2;
  assign c_h_1_28 = c_h_1_24 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3;
  assign c_h_1_29 = c_h_1_21 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_30 = c_h_1_14 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6
      = (mantissa[11:10]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1
      & c_h_1_27 & c_h_1_28 & c_h_1_29;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2
      = ~((mantissa[7:6]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1
      = ~((mantissa[9:8]!=2'b00));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1
      = ~((mantissa[5:4]!=2'b00));
  assign c_h_1_33 = ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1
      & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3
      = (mantissa[3:2]==2'b00) & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1;
  assign c_h_1_34 = c_h_1_33 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3;
  assign c_h_1_35 = c_h_1_30 & ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc
      = (mantissa[1:0]==2'b00) & c_h_1_34 & c_h_1_35;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_nl
      = c_h_1_30 & (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_186_6_sdt_6);
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_1_nl
      = c_h_1_14 & (c_h_1_29 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_90_5_sdt_5))
      & (~ c_h_1_35);
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_292_nl
      = c_h_1_6 & (c_h_1_13 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_42_4_sdt_4))
      & (~((~(c_h_1_21 & (c_h_1_28 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_134_4_sdt_4))))
      & c_h_1_30)) & (c_h_1_34 | (~ c_h_1_35));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_2_nl
      = c_h_1_2 & (c_h_1_5 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_18_3_sdt_3))
      & (~((~(c_h_1_9 & (c_h_1_12 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~((~(c_h_1_17 & (c_h_1_20 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_110_3_sdt_3))
      & (~((~(c_h_1_24 & (c_h_1_27 | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_154_3_sdt_3))))
      & c_h_1_29)))) & c_h_1_30)) & (~((~(c_h_1_33 & (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_206_3_sdt_3)))
      & c_h_1_35));
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_or_2_nl
      = (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_14_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_34_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_58_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_50_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_78_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_106_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_98_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_126_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_118_2_sdt_2))))
      & c_h_1_21)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_150_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_142_2_sdt_2))
      & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_170_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_162_2_sdt_2))))
      & c_h_1_28)))) & c_h_1_29)))) & c_h_1_30)) & (~((~(ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_1
      & (ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_202_2_sdt_1
      | (~ ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_wrs_c_194_2_sdt_2))
      & (~ c_h_1_34))) & c_h_1_35))) | ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc;
  assign ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_nor_nl
      = ~((mantissa[73]) | (~((mantissa[72:71]!=2'b01))) | (((mantissa[69]) | (~((mantissa[68:67]!=2'b01))))
      & c_h_1_2) | ((~((~((mantissa[65]) | (~((mantissa[64:63]!=2'b01))))) & (~(((mantissa[61])
      | (~((mantissa[60:59]!=2'b01)))) & c_h_1_5)))) & c_h_1_6) | ((~((~((mantissa[57])
      | (~((mantissa[56:55]!=2'b01))))) & (~(((mantissa[53]) | (~((mantissa[52:51]!=2'b01))))
      & c_h_1_9)) & (~((~((~((mantissa[49]) | (~((mantissa[48:47]!=2'b01))))) & (~(((mantissa[45])
      | (~((mantissa[44:43]!=2'b01)))) & c_h_1_12)))) & c_h_1_13)))) & c_h_1_14)
      | ((~((~((mantissa[41]) | (~((mantissa[40:39]!=2'b01))))) & (~(((mantissa[37])
      | (~((mantissa[36:35]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[33]) | (~((mantissa[32:31]!=2'b01)))))
      & (~(((mantissa[29]) | (~((mantissa[28:27]!=2'b01)))) & c_h_1_20)))) & c_h_1_21))
      & (~((~((~((mantissa[25]) | (~((mantissa[24:23]!=2'b01))))) & (~(((mantissa[21])
      | (~((mantissa[20:19]!=2'b01)))) & c_h_1_24)) & (~((~((~((mantissa[17]) | (~((mantissa[16:15]!=2'b01)))))
      & (~(((mantissa[13]) | (~((mantissa[12:11]!=2'b01)))) & c_h_1_27)))) & c_h_1_28))))
      & c_h_1_29)))) & c_h_1_30) | ((~((~((mantissa[9]) | (~((mantissa[8:7]!=2'b01)))))
      & (~(((mantissa[5]) | (~((mantissa[4:3]!=2'b01)))) & c_h_1_33)) & (~((mantissa[1])
      & c_h_1_34)))) & c_h_1_35) | ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_291_ssc);
  assign rtn = {c_h_1_35 , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_1_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_292_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_and_2_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_or_2_nl
      , ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_leading_1_leading_sign_74_0_rtn_nor_nl};
endmodule




//------> /opt/cad/catapult/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Single Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)

module BLOCK_1R1W_RBW #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 
  
)( clk,clken,d,q,radr,wadr,we);

  input  clk;
  input  clken;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" *)
  reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block"
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clk ENABLE clken DATA_OUT q ADDRESS radr
  // writeA :: CLOCK clk ENABLE clken DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clk) begin
        if (clken) begin
          radr_reg <= radr;
        end
      end
      always @(posedge clk) begin
        if (clken) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr_reg];
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clk) begin
        if (clken) begin
            ramq <= mem[radr];
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clk) begin
        if (clken) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clk) begin
        if (clken) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clk) begin
        if (clken) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./softmax_sysc.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5a/871028 Production Release
//  HLS Date:       Tue Apr 14 07:55:32 PDT 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Tue Jun  9 14:16:48 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_12_7_67_128_128_67_1_gen
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_12_7_67_128_128_67_1_gen
    (
  clken, q, radr, we, d, wadr, clken_d, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [66:0] q;
  output [6:0] radr;
  output we;
  output [66:0] d;
  output [6:0] wadr;
  input clken_d;
  input [66:0] d_d;
  output [66:0] q_d;
  input [6:0] radr_d;
  input [6:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_run_fsm (
  clk, rst, run_wen, fsm_output, CONFIG_LOOP_C_0_tr0, BATCH_LOOP_C_0_tr0
);
  input clk;
  input rst;
  input run_wen;
  output [6:0] fsm_output;
  reg [6:0] fsm_output;
  input CONFIG_LOOP_C_0_tr0;
  input BATCH_LOOP_C_0_tr0;


  // FSM State Type Declaration for esp_acc_softmax_sysc_softmax_sysc_run_run_fsm_1
  parameter
    run_rlp_C_0 = 3'd0,
    CONFIG_LOOP_C_0 = 3'd1,
    BATCH_LOOP_C_0 = 3'd2,
    run_rlp_C_1 = 3'd3,
    run_rlp_C_2 = 3'd4,
    run_rlp_C_3 = 3'd5,
    PROCESS_DONE_LOOP_C_0 = 3'd6;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : esp_acc_softmax_sysc_softmax_sysc_run_run_fsm_1
    case (state_var)
      CONFIG_LOOP_C_0 : begin
        fsm_output = 7'b0000010;
        if ( CONFIG_LOOP_C_0_tr0 ) begin
          state_var_NS = CONFIG_LOOP_C_0;
        end
        else begin
          state_var_NS = BATCH_LOOP_C_0;
        end
      end
      BATCH_LOOP_C_0 : begin
        fsm_output = 7'b0000100;
        if ( BATCH_LOOP_C_0_tr0 ) begin
          state_var_NS = BATCH_LOOP_C_0;
        end
        else begin
          state_var_NS = run_rlp_C_1;
        end
      end
      run_rlp_C_1 : begin
        fsm_output = 7'b0001000;
        state_var_NS = run_rlp_C_2;
      end
      run_rlp_C_2 : begin
        fsm_output = 7'b0010000;
        state_var_NS = run_rlp_C_3;
      end
      run_rlp_C_3 : begin
        fsm_output = 7'b0100000;
        state_var_NS = PROCESS_DONE_LOOP_C_0;
      end
      PROCESS_DONE_LOOP_C_0 : begin
        fsm_output = 7'b1000000;
        state_var_NS = PROCESS_DONE_LOOP_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 7'b0000001;
        state_var_NS = CONFIG_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( ~ rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_staller
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_staller (
  clk, rst, run_wen, run_wten, dma_read_ctrl_Push_mioi_wen_comp, dma_read_chnl_Pop_mioi_wen_comp,
      dma_write_ctrl_Push_mioi_wen_comp, dma_write_chnl_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output run_wen;
  output run_wten;
  input dma_read_ctrl_Push_mioi_wen_comp;
  input dma_read_chnl_Pop_mioi_wen_comp;
  input dma_write_ctrl_Push_mioi_wen_comp;
  input dma_write_chnl_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg run_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign run_wen = dma_read_ctrl_Push_mioi_wen_comp & dma_read_chnl_Pop_mioi_wen_comp
      & dma_write_ctrl_Push_mioi_wen_comp & dma_write_chnl_Push_mioi_wen_comp;
  assign run_wten = run_wten_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      run_wten_reg <= 1'b0;
    end
    else begin
      run_wten_reg <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_dp
    (
  clk, rst, CALC_SOFTMAX_LOOP_mul_cmp_bawt, CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt, CALC_SOFTMAX_LOOP_mul_cmp_biwt,
      CALC_SOFTMAX_LOOP_mul_cmp_bdwt, CALC_SOFTMAX_LOOP_mul_cmp_z
);
  input clk;
  input rst;
  output CALC_SOFTMAX_LOOP_mul_cmp_bawt;
  output [31:0] CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt;
  input CALC_SOFTMAX_LOOP_mul_cmp_biwt;
  input CALC_SOFTMAX_LOOP_mul_cmp_bdwt;
  input [94:0] CALC_SOFTMAX_LOOP_mul_cmp_z;


  // Interconnect Declarations
  reg [1:0] CALC_SOFTMAX_LOOP_mul_cmp_bcwt;
  wire [2:0] nl_CALC_SOFTMAX_LOOP_mul_cmp_bcwt;
  reg [31:0] CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_2_94_63;
  reg [31:0] CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_1_94_63;
  reg [31:0] CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_94_63;

  wire[1:0] CALC_SOFTMAX_LOOP_acc_1_nl;
  wire[2:0] nl_CALC_SOFTMAX_LOOP_acc_1_nl;
  wire[1:0] CALC_SOFTMAX_LOOP_acc_2_nl;
  wire[2:0] nl_CALC_SOFTMAX_LOOP_acc_2_nl;

  // Interconnect Declarations for Component Instantiations 
  assign CALC_SOFTMAX_LOOP_mul_cmp_bawt = CALC_SOFTMAX_LOOP_mul_cmp_biwt | (CALC_SOFTMAX_LOOP_mul_cmp_bcwt!=2'b00);
  assign CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt = MUX_v_32_4_2((CALC_SOFTMAX_LOOP_mul_cmp_z[94:63]),
      CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_94_63, CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_1_94_63,
      CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_2_94_63, CALC_SOFTMAX_LOOP_mul_cmp_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_mul_cmp_bcwt <= 2'b00;
    end
    else begin
      CALC_SOFTMAX_LOOP_mul_cmp_bcwt <= nl_CALC_SOFTMAX_LOOP_mul_cmp_bcwt[1:0];
    end
  end
  always @(posedge clk) begin
    if ( CALC_SOFTMAX_LOOP_mul_cmp_biwt ) begin
      CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_94_63 <= CALC_SOFTMAX_LOOP_mul_cmp_z[94:63];
      CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_1_94_63 <= CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_94_63;
      CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_2_94_63 <= CALC_SOFTMAX_LOOP_mul_cmp_z_bfwt_1_94_63;
    end
  end
  assign nl_CALC_SOFTMAX_LOOP_acc_1_nl = conv_u2u_1_2(CALC_SOFTMAX_LOOP_mul_cmp_biwt)
      + conv_u2u_1_2(~ CALC_SOFTMAX_LOOP_mul_cmp_bdwt);
  assign CALC_SOFTMAX_LOOP_acc_1_nl = nl_CALC_SOFTMAX_LOOP_acc_1_nl[1:0];
  assign nl_CALC_SOFTMAX_LOOP_acc_2_nl = CALC_SOFTMAX_LOOP_mul_cmp_bcwt + 2'b11;
  assign CALC_SOFTMAX_LOOP_acc_2_nl = nl_CALC_SOFTMAX_LOOP_acc_2_nl[1:0];
  assign nl_CALC_SOFTMAX_LOOP_mul_cmp_bcwt  = CALC_SOFTMAX_LOOP_acc_1_nl + CALC_SOFTMAX_LOOP_acc_2_nl;

  function automatic [31:0] MUX_v_32_4_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [31:0] input_3;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_32_4_2 = result;
  end
  endfunction


  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_ctrl
    (
  clk, rst, run_wen, run_wten, CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg, CALC_SOFTMAX_LOOP_mul_cmp_iswt2,
      CALC_SOFTMAX_LOOP_mul_cmp_biwt, CALC_SOFTMAX_LOOP_mul_cmp_bdwt
);
  input clk;
  input rst;
  input run_wen;
  input run_wten;
  input CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg;
  input CALC_SOFTMAX_LOOP_mul_cmp_iswt2;
  output CALC_SOFTMAX_LOOP_mul_cmp_biwt;
  output CALC_SOFTMAX_LOOP_mul_cmp_bdwt;


  // Interconnect Declarations
  reg CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt1;
  reg CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt0;
  reg [1:0] CALC_SOFTMAX_LOOP_mul_cmp_icwt;
  wire [2:0] nl_CALC_SOFTMAX_LOOP_mul_cmp_icwt;

  wire[1:0] CALC_SOFTMAX_LOOP_acc_2_nl;
  wire[2:0] nl_CALC_SOFTMAX_LOOP_acc_2_nl;
  wire[1:0] CALC_SOFTMAX_LOOP_acc_3_nl;
  wire[2:0] nl_CALC_SOFTMAX_LOOP_acc_3_nl;

  // Interconnect Declarations for Component Instantiations 
  assign CALC_SOFTMAX_LOOP_mul_cmp_bdwt = CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg &
      run_wen;
  assign CALC_SOFTMAX_LOOP_mul_cmp_biwt = CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt0
      | (CALC_SOFTMAX_LOOP_mul_cmp_icwt!=2'b00);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt1 <= 1'b0;
      CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt0 <= 1'b0;
      CALC_SOFTMAX_LOOP_mul_cmp_icwt <= 2'b00;
    end
    else begin
      CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt1 <= (~ run_wten) &
          CALC_SOFTMAX_LOOP_mul_cmp_iswt2;
      CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt0 <= CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt1;
      CALC_SOFTMAX_LOOP_mul_cmp_icwt <= nl_CALC_SOFTMAX_LOOP_mul_cmp_icwt[1:0];
    end
  end
  assign nl_CALC_SOFTMAX_LOOP_acc_2_nl = conv_u2u_1_2(CALC_SOFTMAX_LOOP_mul_cmp_ALC_SOFTMAX_LOOP_mul_cmp_pdswt0)
      + conv_u2u_1_2(~ CALC_SOFTMAX_LOOP_mul_cmp_biwt);
  assign CALC_SOFTMAX_LOOP_acc_2_nl = nl_CALC_SOFTMAX_LOOP_acc_2_nl[1:0];
  assign nl_CALC_SOFTMAX_LOOP_acc_3_nl = CALC_SOFTMAX_LOOP_mul_cmp_icwt + 2'b11;
  assign CALC_SOFTMAX_LOOP_acc_3_nl = nl_CALC_SOFTMAX_LOOP_acc_3_nl[1:0];
  assign nl_CALC_SOFTMAX_LOOP_mul_cmp_icwt  = CALC_SOFTMAX_LOOP_acc_2_nl + CALC_SOFTMAX_LOOP_acc_3_nl;

  function automatic [1:0] conv_u2u_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_2 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_dp
    (
  clk, rst, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2
);
  input clk;
  input rst;
  input [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt;
  output [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2;


  // Interconnect Declarations
  reg ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt;
  reg ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt_1;
  reg [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt
      | ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt
      = MUX_v_67_2_2(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_bfwt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt_1);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt
          <= 1'b0;
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt_1
          <= 1'b0;
    end
    else begin
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt
          <= ~((~(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt
          | ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt))
          | ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt);
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt_1
          <= ~((~(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bcwt_1
          | ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1))
          | ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2);
    end
  end
  always @(posedge clk) begin
    if ( ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1
        ) begin
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_bfwt
          <= ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d;
    end
  end

  function automatic [66:0] MUX_v_67_2_2;
    input [66:0] input_0;
    input [66:0] input_1;
    input [0:0] sel;
    reg [66:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_67_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_ctrl
    (
  run_wen, run_wten, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_run_sct,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_run_sct_pff,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff
);
  input run_wen;
  input run_wten;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_run_sct;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_run_sct_pff;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg
      & run_wen;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt
      = (~ run_wten) & ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1
      & run_wen;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1
      = (~ run_wten) & ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_run_sct_pff
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff
      & run_wen;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_run_sct
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff
      & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp
    (
  clk, rst, dma_write_chnl_Push_mioi_oswt_unreg, dma_write_chnl_Push_mioi_bawt, dma_write_chnl_Push_mioi_wen_comp,
      dma_write_chnl_Push_mioi_biwt, dma_write_chnl_Push_mioi_bdwt
);
  input clk;
  input rst;
  input dma_write_chnl_Push_mioi_oswt_unreg;
  output dma_write_chnl_Push_mioi_bawt;
  output dma_write_chnl_Push_mioi_wen_comp;
  input dma_write_chnl_Push_mioi_biwt;
  input dma_write_chnl_Push_mioi_bdwt;


  // Interconnect Declarations
  reg dma_write_chnl_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_write_chnl_Push_mioi_bawt = dma_write_chnl_Push_mioi_biwt | dma_write_chnl_Push_mioi_bcwt;
  assign dma_write_chnl_Push_mioi_wen_comp = (~ dma_write_chnl_Push_mioi_oswt_unreg)
      | dma_write_chnl_Push_mioi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_chnl_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_write_chnl_Push_mioi_bcwt <= ~((~(dma_write_chnl_Push_mioi_bcwt | dma_write_chnl_Push_mioi_biwt))
          | dma_write_chnl_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl
    (
  clk, rst, run_wen, run_wten, dma_write_chnl_Push_mioi_oswt_unreg, dma_write_chnl_Push_mioi_iswt0,
      dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct, dma_write_chnl_Push_mioi_biwt,
      dma_write_chnl_Push_mioi_bdwt, dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct,
      dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld, dma_write_chnl_Push_mioi_iswt0_pff
);
  input clk;
  input rst;
  input run_wen;
  input run_wten;
  input dma_write_chnl_Push_mioi_oswt_unreg;
  input dma_write_chnl_Push_mioi_iswt0;
  input dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct;
  output dma_write_chnl_Push_mioi_biwt;
  output dma_write_chnl_Push_mioi_bdwt;
  output dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct;
  input dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld;
  input dma_write_chnl_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire dma_write_chnl_Push_mioi_ogwt;
  reg dma_write_chnl_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_write_chnl_Push_mioi_bdwt = dma_write_chnl_Push_mioi_oswt_unreg & run_wen;
  assign dma_write_chnl_Push_mioi_biwt = dma_write_chnl_Push_mioi_ogwt & dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld;
  assign dma_write_chnl_Push_mioi_ogwt = ((~ run_wten) & dma_write_chnl_Push_mioi_iswt0)
      | dma_write_chnl_Push_mioi_icwt;
  assign dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct = dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct
      & run_wen & dma_write_chnl_Push_mioi_iswt0_pff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_chnl_Push_mioi_icwt <= 1'b0;
    end
    else begin
      dma_write_chnl_Push_mioi_icwt <= dma_write_chnl_Push_mioi_ogwt & (~ dma_write_chnl_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp
    (
  clk, rst, dma_write_ctrl_Push_mioi_oswt_unreg, dma_write_ctrl_Push_mioi_bawt, dma_write_ctrl_Push_mioi_wen_comp,
      dma_write_ctrl_Push_mioi_biwt, dma_write_ctrl_Push_mioi_bdwt
);
  input clk;
  input rst;
  input dma_write_ctrl_Push_mioi_oswt_unreg;
  output dma_write_ctrl_Push_mioi_bawt;
  output dma_write_ctrl_Push_mioi_wen_comp;
  input dma_write_ctrl_Push_mioi_biwt;
  input dma_write_ctrl_Push_mioi_bdwt;


  // Interconnect Declarations
  reg dma_write_ctrl_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_write_ctrl_Push_mioi_bawt = dma_write_ctrl_Push_mioi_biwt | dma_write_ctrl_Push_mioi_bcwt;
  assign dma_write_ctrl_Push_mioi_wen_comp = (~ dma_write_ctrl_Push_mioi_oswt_unreg)
      | dma_write_ctrl_Push_mioi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_ctrl_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_write_ctrl_Push_mioi_bcwt <= ~((~(dma_write_ctrl_Push_mioi_bcwt | dma_write_ctrl_Push_mioi_biwt))
          | dma_write_ctrl_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl
    (
  clk, rst, run_wen, run_wten, dma_write_ctrl_Push_mioi_oswt_unreg, dma_write_ctrl_Push_mioi_iswt0,
      dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct, dma_write_ctrl_Push_mioi_biwt,
      dma_write_ctrl_Push_mioi_bdwt, dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct,
      dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld, dma_write_ctrl_Push_mioi_iswt0_pff
);
  input clk;
  input rst;
  input run_wen;
  input run_wten;
  input dma_write_ctrl_Push_mioi_oswt_unreg;
  input dma_write_ctrl_Push_mioi_iswt0;
  input dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct;
  output dma_write_ctrl_Push_mioi_biwt;
  output dma_write_ctrl_Push_mioi_bdwt;
  output dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct;
  input dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  input dma_write_ctrl_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire dma_write_ctrl_Push_mioi_ogwt;
  reg dma_write_ctrl_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_write_ctrl_Push_mioi_bdwt = dma_write_ctrl_Push_mioi_oswt_unreg & run_wen;
  assign dma_write_ctrl_Push_mioi_biwt = dma_write_ctrl_Push_mioi_ogwt & dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  assign dma_write_ctrl_Push_mioi_ogwt = ((~ run_wten) & dma_write_ctrl_Push_mioi_iswt0)
      | dma_write_ctrl_Push_mioi_icwt;
  assign dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct = dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct
      & run_wen & dma_write_ctrl_Push_mioi_iswt0_pff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_write_ctrl_Push_mioi_icwt <= 1'b0;
    end
    else begin
      dma_write_ctrl_Push_mioi_icwt <= dma_write_ctrl_Push_mioi_ogwt & (~ dma_write_ctrl_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp
    (
  clk, rst, dma_read_chnl_Pop_mioi_oswt_unreg, dma_read_chnl_Pop_mioi_bawt, dma_read_chnl_Pop_mioi_wen_comp,
      dma_read_chnl_Pop_mioi_return_rsc_z_mxwt, dma_read_chnl_Pop_mioi_return_rsc_z,
      dma_read_chnl_Pop_mioi_biwt, dma_read_chnl_Pop_mioi_bdwt
);
  input clk;
  input rst;
  input dma_read_chnl_Pop_mioi_oswt_unreg;
  output dma_read_chnl_Pop_mioi_bawt;
  output dma_read_chnl_Pop_mioi_wen_comp;
  output [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt;
  input [63:0] dma_read_chnl_Pop_mioi_return_rsc_z;
  input dma_read_chnl_Pop_mioi_biwt;
  input dma_read_chnl_Pop_mioi_bdwt;


  // Interconnect Declarations
  reg dma_read_chnl_Pop_mioi_bcwt;
  reg [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_bfwt_31_0;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_chnl_Pop_mioi_bawt = dma_read_chnl_Pop_mioi_biwt | dma_read_chnl_Pop_mioi_bcwt;
  assign dma_read_chnl_Pop_mioi_wen_comp = (~ dma_read_chnl_Pop_mioi_oswt_unreg)
      | dma_read_chnl_Pop_mioi_bawt;
  assign dma_read_chnl_Pop_mioi_return_rsc_z_mxwt = MUX_v_32_2_2((dma_read_chnl_Pop_mioi_return_rsc_z[31:0]),
      dma_read_chnl_Pop_mioi_return_rsc_z_bfwt_31_0, dma_read_chnl_Pop_mioi_bcwt);
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_chnl_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_read_chnl_Pop_mioi_bcwt <= ~((~(dma_read_chnl_Pop_mioi_bcwt | dma_read_chnl_Pop_mioi_biwt))
          | dma_read_chnl_Pop_mioi_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( dma_read_chnl_Pop_mioi_biwt ) begin
      dma_read_chnl_Pop_mioi_return_rsc_z_bfwt_31_0 <= dma_read_chnl_Pop_mioi_return_rsc_z[31:0];
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl
    (
  clk, rst, run_wen, run_wten, dma_read_chnl_Pop_mioi_oswt_unreg, dma_read_chnl_Pop_mioi_iswt0,
      dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_psct, dma_read_chnl_Pop_mioi_biwt,
      dma_read_chnl_Pop_mioi_bdwt, dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct,
      dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld, dma_read_chnl_Pop_mioi_iswt0_pff
);
  input clk;
  input rst;
  input run_wen;
  input run_wten;
  input dma_read_chnl_Pop_mioi_oswt_unreg;
  input dma_read_chnl_Pop_mioi_iswt0;
  input dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_psct;
  output dma_read_chnl_Pop_mioi_biwt;
  output dma_read_chnl_Pop_mioi_bdwt;
  output dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct;
  input dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld;
  input dma_read_chnl_Pop_mioi_iswt0_pff;


  // Interconnect Declarations
  wire dma_read_chnl_Pop_mioi_ogwt;
  reg dma_read_chnl_Pop_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_chnl_Pop_mioi_bdwt = dma_read_chnl_Pop_mioi_oswt_unreg & run_wen;
  assign dma_read_chnl_Pop_mioi_biwt = dma_read_chnl_Pop_mioi_ogwt & dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld;
  assign dma_read_chnl_Pop_mioi_ogwt = ((~ run_wten) & dma_read_chnl_Pop_mioi_iswt0)
      | dma_read_chnl_Pop_mioi_icwt;
  assign dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct = dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_psct
      & run_wen & dma_read_chnl_Pop_mioi_iswt0_pff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_chnl_Pop_mioi_icwt <= 1'b0;
    end
    else begin
      dma_read_chnl_Pop_mioi_icwt <= dma_read_chnl_Pop_mioi_ogwt & (~ dma_read_chnl_Pop_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp
    (
  clk, rst, dma_read_ctrl_Push_mioi_oswt_unreg, dma_read_ctrl_Push_mioi_bawt, dma_read_ctrl_Push_mioi_wen_comp,
      dma_read_ctrl_Push_mioi_biwt, dma_read_ctrl_Push_mioi_bdwt
);
  input clk;
  input rst;
  input dma_read_ctrl_Push_mioi_oswt_unreg;
  output dma_read_ctrl_Push_mioi_bawt;
  output dma_read_ctrl_Push_mioi_wen_comp;
  input dma_read_ctrl_Push_mioi_biwt;
  input dma_read_ctrl_Push_mioi_bdwt;


  // Interconnect Declarations
  reg dma_read_ctrl_Push_mioi_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_ctrl_Push_mioi_bawt = dma_read_ctrl_Push_mioi_biwt | dma_read_ctrl_Push_mioi_bcwt;
  assign dma_read_ctrl_Push_mioi_wen_comp = (~ dma_read_ctrl_Push_mioi_oswt_unreg)
      | dma_read_ctrl_Push_mioi_bawt;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      dma_read_ctrl_Push_mioi_bcwt <= ~((~(dma_read_ctrl_Push_mioi_bcwt | dma_read_ctrl_Push_mioi_biwt))
          | dma_read_ctrl_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl
    (
  clk, rst, run_wen, dma_read_ctrl_Push_mioi_oswt_unreg, dma_read_ctrl_Push_mioi_iswt0,
      run_wten, dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct, dma_read_ctrl_Push_mioi_biwt,
      dma_read_ctrl_Push_mioi_bdwt, dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct,
      dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld, dma_read_ctrl_Push_mioi_iswt0_pff
);
  input clk;
  input rst;
  input run_wen;
  input dma_read_ctrl_Push_mioi_oswt_unreg;
  input dma_read_ctrl_Push_mioi_iswt0;
  input run_wten;
  input dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct;
  output dma_read_ctrl_Push_mioi_biwt;
  output dma_read_ctrl_Push_mioi_bdwt;
  output dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct;
  input dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  input dma_read_ctrl_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire dma_read_ctrl_Push_mioi_ogwt;
  reg dma_read_ctrl_Push_mioi_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign dma_read_ctrl_Push_mioi_bdwt = dma_read_ctrl_Push_mioi_oswt_unreg & run_wen;
  assign dma_read_ctrl_Push_mioi_biwt = dma_read_ctrl_Push_mioi_ogwt & dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld;
  assign dma_read_ctrl_Push_mioi_ogwt = ((~ run_wten) & dma_read_ctrl_Push_mioi_iswt0)
      | dma_read_ctrl_Push_mioi_icwt;
  assign dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct = dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct
      & run_wen & dma_read_ctrl_Push_mioi_iswt0_pff;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_Push_mioi_icwt <= 1'b0;
    end
    else begin
      dma_read_ctrl_Push_mioi_icwt <= dma_read_ctrl_Push_mioi_ogwt & (~ dma_read_ctrl_Push_mioi_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp (
  clk, rst, run_wen, run_wten, CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg, CALC_SOFTMAX_LOOP_mul_cmp_bawt,
      CALC_SOFTMAX_LOOP_mul_cmp_iswt2, CALC_SOFTMAX_LOOP_mul_cmp_a_run, CALC_SOFTMAX_LOOP_mul_cmp_b_run,
      CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt
);
  input clk;
  input rst;
  input run_wen;
  input run_wten;
  input CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg;
  output CALC_SOFTMAX_LOOP_mul_cmp_bawt;
  input CALC_SOFTMAX_LOOP_mul_cmp_iswt2;
  input [66:0] CALC_SOFTMAX_LOOP_mul_cmp_a_run;
  input [93:0] CALC_SOFTMAX_LOOP_mul_cmp_b_run;
  output [31:0] CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt;


  // Interconnect Declarations
  wire CALC_SOFTMAX_LOOP_mul_cmp_biwt;
  wire CALC_SOFTMAX_LOOP_mul_cmp_bdwt;
  wire [94:0] CALC_SOFTMAX_LOOP_mul_cmp_z;
  wire [31:0] CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_mgc_mul_pipe #(.width_a(32'sd67),
  .signd_a(32'sd0),
  .width_b(32'sd94),
  .signd_b(32'sd0),
  .width_z(32'sd95),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) CALC_SOFTMAX_LOOP_mul_cmp (
      .a(CALC_SOFTMAX_LOOP_mul_cmp_a_run),
      .b(CALC_SOFTMAX_LOOP_mul_cmp_b_run),
      .clk(clk),
      .en(1'b1),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(CALC_SOFTMAX_LOOP_mul_cmp_z)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_ctrl
      softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg(CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg),
      .CALC_SOFTMAX_LOOP_mul_cmp_iswt2(CALC_SOFTMAX_LOOP_mul_cmp_iswt2),
      .CALC_SOFTMAX_LOOP_mul_cmp_biwt(CALC_SOFTMAX_LOOP_mul_cmp_biwt),
      .CALC_SOFTMAX_LOOP_mul_cmp_bdwt(CALC_SOFTMAX_LOOP_mul_cmp_bdwt)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_dp
      softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp_mgc_mul_pipe_67_0_94_0_95_1_1_0_0_3_1_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .CALC_SOFTMAX_LOOP_mul_cmp_bawt(CALC_SOFTMAX_LOOP_mul_cmp_bawt),
      .CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt(CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt_pconst),
      .CALC_SOFTMAX_LOOP_mul_cmp_biwt(CALC_SOFTMAX_LOOP_mul_cmp_biwt),
      .CALC_SOFTMAX_LOOP_mul_cmp_bdwt(CALC_SOFTMAX_LOOP_mul_cmp_bdwt),
      .CALC_SOFTMAX_LOOP_mul_cmp_z(CALC_SOFTMAX_LOOP_mul_cmp_z)
    );
  assign CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt = CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1
    (
  clk, rst, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      run_wen, run_wten, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff
);
  input clk;
  input rst;
  input [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  input run_wen;
  input run_wten;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1;
  output [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff;
  input ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff;


  // Interconnect Declarations
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_run_sct;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_ctrl
      softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_run_sct(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_run_sct),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_run_sct_pff(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_run_sct_iff),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_dp
      softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_biwt_1),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bdwt_2)
    );
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_run_sct_iff;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_run_sct;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_dma_write_chnl_Push_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_dma_write_chnl_Push_mioi (
  clk, rst, dma_write_chnl_val, dma_write_chnl_rdy, dma_write_chnl_msg, run_wen,
      run_wten, dma_write_chnl_Push_mioi_m_rsc_dat, dma_write_chnl_Push_mioi_oswt_unreg,
      dma_write_chnl_Push_mioi_bawt, dma_write_chnl_Push_mioi_iswt0, dma_write_chnl_Push_mioi_wen_comp,
      dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct, dma_write_chnl_Push_mioi_iswt0_pff
);
  input clk;
  input rst;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;
  input run_wen;
  input run_wten;
  input [63:0] dma_write_chnl_Push_mioi_m_rsc_dat;
  input dma_write_chnl_Push_mioi_oswt_unreg;
  output dma_write_chnl_Push_mioi_bawt;
  input dma_write_chnl_Push_mioi_iswt0;
  output dma_write_chnl_Push_mioi_wen_comp;
  input dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct;
  input dma_write_chnl_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire dma_write_chnl_Push_mioi_biwt;
  wire dma_write_chnl_Push_mioi_bdwt;
  wire dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct;
  wire dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  wire [63:0] nl_dma_write_chnl_Push_mioi_m_rsc_dat;
  assign nl_dma_write_chnl_Push_mioi_m_rsc_dat = {32'b11011110101011011011111011101111
      , (dma_write_chnl_Push_mioi_m_rsc_dat[31:0])};
  esp_acc_softmax_sysc_Connections_OutBlocking_dma_data_t_Connections_SYN_PORT_Push
      dma_write_chnl_Push_mioi (
      .this_val(dma_write_chnl_val),
      .this_rdy(dma_write_chnl_rdy),
      .this_msg(dma_write_chnl_msg),
      .m_rsc_dat(nl_dma_write_chnl_Push_mioi_m_rsc_dat[63:0]),
      .ccs_ccore_start_rsc_dat(dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .ccs_ccore_done_sync_vld(dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl
      softmax_sysc_run_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .dma_write_chnl_Push_mioi_oswt_unreg(dma_write_chnl_Push_mioi_oswt_unreg),
      .dma_write_chnl_Push_mioi_iswt0(dma_write_chnl_Push_mioi_iswt0),
      .dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct(dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct),
      .dma_write_chnl_Push_mioi_biwt(dma_write_chnl_Push_mioi_biwt),
      .dma_write_chnl_Push_mioi_bdwt(dma_write_chnl_Push_mioi_bdwt),
      .dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct(dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld(dma_write_chnl_Push_mioi_ccs_ccore_done_sync_vld),
      .dma_write_chnl_Push_mioi_iswt0_pff(dma_write_chnl_Push_mioi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp
      softmax_sysc_run_dma_write_chnl_Push_mioi_dma_write_chnl_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_chnl_Push_mioi_oswt_unreg(dma_write_chnl_Push_mioi_oswt_unreg),
      .dma_write_chnl_Push_mioi_bawt(dma_write_chnl_Push_mioi_bawt),
      .dma_write_chnl_Push_mioi_wen_comp(dma_write_chnl_Push_mioi_wen_comp),
      .dma_write_chnl_Push_mioi_biwt(dma_write_chnl_Push_mioi_biwt),
      .dma_write_chnl_Push_mioi_bdwt(dma_write_chnl_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_dma_write_ctrl_Push_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_dma_write_ctrl_Push_mioi (
  clk, rst, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg, run_wen,
      run_wten, dma_write_ctrl_Push_mioi_m_index_rsc_dat, dma_write_ctrl_Push_mioi_oswt_unreg,
      dma_write_ctrl_Push_mioi_bawt, dma_write_ctrl_Push_mioi_iswt0, dma_write_ctrl_Push_mioi_wen_comp,
      dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct, dma_write_ctrl_Push_mioi_iswt0_pff
);
  input clk;
  input rst;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  input run_wen;
  input run_wten;
  input [31:0] dma_write_ctrl_Push_mioi_m_index_rsc_dat;
  input dma_write_ctrl_Push_mioi_oswt_unreg;
  output dma_write_ctrl_Push_mioi_bawt;
  input dma_write_ctrl_Push_mioi_iswt0;
  output dma_write_ctrl_Push_mioi_wen_comp;
  input dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct;
  input dma_write_ctrl_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire dma_write_ctrl_Push_mioi_biwt;
  wire dma_write_ctrl_Push_mioi_bdwt;
  wire dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct;
  wire dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_dma_write_ctrl_Push_mioi_m_index_rsc_dat;
  assign nl_dma_write_ctrl_Push_mioi_m_index_rsc_dat = {(dma_write_ctrl_Push_mioi_m_index_rsc_dat[31:7])
      , 7'b0000000};
  esp_acc_softmax_sysc_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push
      dma_write_ctrl_Push_mioi (
      .this_val(dma_write_ctrl_val),
      .this_rdy(dma_write_ctrl_rdy),
      .this_msg(dma_write_ctrl_msg),
      .m_index_rsc_dat(nl_dma_write_ctrl_Push_mioi_m_index_rsc_dat[31:0]),
      .ccs_ccore_start_rsc_dat(dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .ccs_ccore_done_sync_vld(dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl
      softmax_sysc_run_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .dma_write_ctrl_Push_mioi_oswt_unreg(dma_write_ctrl_Push_mioi_oswt_unreg),
      .dma_write_ctrl_Push_mioi_iswt0(dma_write_ctrl_Push_mioi_iswt0),
      .dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct(dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct),
      .dma_write_ctrl_Push_mioi_biwt(dma_write_ctrl_Push_mioi_biwt),
      .dma_write_ctrl_Push_mioi_bdwt(dma_write_ctrl_Push_mioi_bdwt),
      .dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct(dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld(dma_write_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .dma_write_ctrl_Push_mioi_iswt0_pff(dma_write_ctrl_Push_mioi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp
      softmax_sysc_run_dma_write_ctrl_Push_mioi_dma_write_ctrl_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_ctrl_Push_mioi_oswt_unreg(dma_write_ctrl_Push_mioi_oswt_unreg),
      .dma_write_ctrl_Push_mioi_bawt(dma_write_ctrl_Push_mioi_bawt),
      .dma_write_ctrl_Push_mioi_wen_comp(dma_write_ctrl_Push_mioi_wen_comp),
      .dma_write_ctrl_Push_mioi_biwt(dma_write_ctrl_Push_mioi_biwt),
      .dma_write_ctrl_Push_mioi_bdwt(dma_write_ctrl_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_dma_read_chnl_Pop_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_dma_read_chnl_Pop_mioi (
  clk, rst, dma_read_chnl_val, dma_read_chnl_rdy, dma_read_chnl_msg, run_wen, run_wten,
      dma_read_chnl_Pop_mioi_oswt_unreg, dma_read_chnl_Pop_mioi_bawt, dma_read_chnl_Pop_mioi_iswt0,
      dma_read_chnl_Pop_mioi_wen_comp, dma_read_chnl_Pop_mioi_return_rsc_z_mxwt,
      dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_psct, dma_read_chnl_Pop_mioi_iswt0_pff
);
  input clk;
  input rst;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  input run_wen;
  input run_wten;
  input dma_read_chnl_Pop_mioi_oswt_unreg;
  output dma_read_chnl_Pop_mioi_bawt;
  input dma_read_chnl_Pop_mioi_iswt0;
  output dma_read_chnl_Pop_mioi_wen_comp;
  output [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt;
  input dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_psct;
  input dma_read_chnl_Pop_mioi_iswt0_pff;


  // Interconnect Declarations
  wire [63:0] dma_read_chnl_Pop_mioi_return_rsc_z;
  wire dma_read_chnl_Pop_mioi_biwt;
  wire dma_read_chnl_Pop_mioi_bdwt;
  wire dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct;
  wire dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld;
  wire [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  esp_acc_softmax_sysc_Connections_InBlocking_dma_data_t_Connections_SYN_PORT_Pop
      dma_read_chnl_Pop_mioi (
      .this_val(dma_read_chnl_val),
      .this_rdy(dma_read_chnl_rdy),
      .this_msg(dma_read_chnl_msg),
      .return_rsc_z(dma_read_chnl_Pop_mioi_return_rsc_z),
      .ccs_ccore_start_rsc_dat(dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .ccs_ccore_done_sync_vld(dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl
      softmax_sysc_run_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .dma_read_chnl_Pop_mioi_oswt_unreg(dma_read_chnl_Pop_mioi_oswt_unreg),
      .dma_read_chnl_Pop_mioi_iswt0(dma_read_chnl_Pop_mioi_iswt0),
      .dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_psct(dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_psct),
      .dma_read_chnl_Pop_mioi_biwt(dma_read_chnl_Pop_mioi_biwt),
      .dma_read_chnl_Pop_mioi_bdwt(dma_read_chnl_Pop_mioi_bdwt),
      .dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct(dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld(dma_read_chnl_Pop_mioi_ccs_ccore_done_sync_vld),
      .dma_read_chnl_Pop_mioi_iswt0_pff(dma_read_chnl_Pop_mioi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp
      softmax_sysc_run_dma_read_chnl_Pop_mioi_dma_read_chnl_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_chnl_Pop_mioi_oswt_unreg(dma_read_chnl_Pop_mioi_oswt_unreg),
      .dma_read_chnl_Pop_mioi_bawt(dma_read_chnl_Pop_mioi_bawt),
      .dma_read_chnl_Pop_mioi_wen_comp(dma_read_chnl_Pop_mioi_wen_comp),
      .dma_read_chnl_Pop_mioi_return_rsc_z_mxwt(dma_read_chnl_Pop_mioi_return_rsc_z_mxwt_pconst),
      .dma_read_chnl_Pop_mioi_return_rsc_z(dma_read_chnl_Pop_mioi_return_rsc_z),
      .dma_read_chnl_Pop_mioi_biwt(dma_read_chnl_Pop_mioi_biwt),
      .dma_read_chnl_Pop_mioi_bdwt(dma_read_chnl_Pop_mioi_bdwt)
    );
  assign dma_read_chnl_Pop_mioi_return_rsc_z_mxwt = dma_read_chnl_Pop_mioi_return_rsc_z_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run_dma_read_ctrl_Push_mioi
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run_dma_read_ctrl_Push_mioi (
  clk, rst, dma_read_ctrl_val, dma_read_ctrl_rdy, dma_read_ctrl_msg, run_wen, dma_read_ctrl_Push_mioi_m_index_rsc_dat,
      dma_read_ctrl_Push_mioi_oswt_unreg, dma_read_ctrl_Push_mioi_bawt, dma_read_ctrl_Push_mioi_iswt0,
      run_wten, dma_read_ctrl_Push_mioi_wen_comp, dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct,
      dma_read_ctrl_Push_mioi_iswt0_pff
);
  input clk;
  input rst;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  input run_wen;
  input [31:0] dma_read_ctrl_Push_mioi_m_index_rsc_dat;
  input dma_read_ctrl_Push_mioi_oswt_unreg;
  output dma_read_ctrl_Push_mioi_bawt;
  input dma_read_ctrl_Push_mioi_iswt0;
  input run_wten;
  output dma_read_ctrl_Push_mioi_wen_comp;
  input dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct;
  input dma_read_ctrl_Push_mioi_iswt0_pff;


  // Interconnect Declarations
  wire dma_read_ctrl_Push_mioi_biwt;
  wire dma_read_ctrl_Push_mioi_bdwt;
  wire dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct;
  wire dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_dma_read_ctrl_Push_mioi_m_index_rsc_dat;
  assign nl_dma_read_ctrl_Push_mioi_m_index_rsc_dat = {21'b000000000000000000000
      , (dma_read_ctrl_Push_mioi_m_index_rsc_dat[10:7]) , 7'b0000000};
  esp_acc_softmax_sysc_Connections_OutBlocking_dma_info_t_Connections_SYN_PORT_Push
      dma_read_ctrl_Push_mioi (
      .this_val(dma_read_ctrl_val),
      .this_rdy(dma_read_ctrl_rdy),
      .this_msg(dma_read_ctrl_msg),
      .m_index_rsc_dat(nl_dma_read_ctrl_Push_mioi_m_index_rsc_dat[31:0]),
      .ccs_ccore_start_rsc_dat(dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .ccs_ccore_done_sync_vld(dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(clk),
      .ccs_MIO_srst(rst)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl
      softmax_sysc_run_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_ctrl_inst
      (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .dma_read_ctrl_Push_mioi_oswt_unreg(dma_read_ctrl_Push_mioi_oswt_unreg),
      .dma_read_ctrl_Push_mioi_iswt0(dma_read_ctrl_Push_mioi_iswt0),
      .run_wten(run_wten),
      .dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct(dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct),
      .dma_read_ctrl_Push_mioi_biwt(dma_read_ctrl_Push_mioi_biwt),
      .dma_read_ctrl_Push_mioi_bdwt(dma_read_ctrl_Push_mioi_bdwt),
      .dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct(dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_sct),
      .dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld(dma_read_ctrl_Push_mioi_ccs_ccore_done_sync_vld),
      .dma_read_ctrl_Push_mioi_iswt0_pff(dma_read_ctrl_Push_mioi_iswt0_pff)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp
      softmax_sysc_run_dma_read_ctrl_Push_mioi_dma_read_ctrl_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_ctrl_Push_mioi_oswt_unreg(dma_read_ctrl_Push_mioi_oswt_unreg),
      .dma_read_ctrl_Push_mioi_bawt(dma_read_ctrl_Push_mioi_bawt),
      .dma_read_ctrl_Push_mioi_wen_comp(dma_read_ctrl_Push_mioi_wen_comp),
      .dma_read_ctrl_Push_mioi_biwt(dma_read_ctrl_Push_mioi_biwt),
      .dma_read_ctrl_Push_mioi_bdwt(dma_read_ctrl_Push_mioi_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    esp_acc_softmax_sysc_softmax_sysc_run
// ------------------------------------------------------------------


module esp_acc_softmax_sysc_softmax_sysc_run (
  clk, rst, conf_info, conf_done, acc_done, dma_read_ctrl_val, dma_read_ctrl_rdy,
      dma_read_ctrl_msg, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg,
      dma_read_chnl_val, dma_read_chnl_rdy, dma_read_chnl_msg, dma_write_chnl_val,
      dma_write_chnl_rdy, dma_write_chnl_msg, ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff
);
  input clk;
  input rst;
  input [31:0] conf_info;
  input conf_done;
  output acc_done;
  reg acc_done;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;
  output [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d;
  input [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d;
  output [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d;
  output [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  output ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire dma_read_ctrl_Push_mioi_bawt;
  reg dma_read_ctrl_Push_mioi_iswt0;
  wire run_wten;
  wire dma_read_ctrl_Push_mioi_wen_comp;
  reg dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct;
  wire dma_read_chnl_Pop_mioi_bawt;
  reg dma_read_chnl_Pop_mioi_iswt0;
  wire dma_read_chnl_Pop_mioi_wen_comp;
  wire [31:0] dma_read_chnl_Pop_mioi_return_rsc_z_mxwt;
  reg dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_psct;
  wire dma_write_ctrl_Push_mioi_bawt;
  reg dma_write_ctrl_Push_mioi_iswt0;
  wire dma_write_ctrl_Push_mioi_wen_comp;
  reg dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct;
  wire dma_write_chnl_Push_mioi_bawt;
  wire dma_write_chnl_Push_mioi_wen_comp;
  reg dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt;
  wire CALC_SOFTMAX_LOOP_mul_cmp_bawt;
  wire [31:0] CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt;
  reg [3:0] dma_read_ctrl_Push_mioi_m_index_rsc_dat_10_7;
  reg [24:0] dma_write_ctrl_Push_mioi_m_index_rsc_dat_31_7;
  reg [31:0] dma_write_chnl_Push_mioi_m_rsc_dat_31_0;
  wire [6:0] fsm_output;
  wire BATCH_LOOP_nor_8_tmp;
  wire [7:0] SUM_EXP_LOOP_acc_2_tmp;
  wire [8:0] nl_SUM_EXP_LOOP_acc_2_tmp;
  wire [7:0] CALC_EXP_LOOP_acc_1_tmp;
  wire [8:0] nl_CALC_EXP_LOOP_acc_1_tmp;
  wire [7:0] LOAD_LOOP_acc_2_tmp;
  wire [8:0] nl_LOAD_LOOP_acc_2_tmp;
  wire [4:0] BATCH_LOOP_acc_3_tmp;
  wire [5:0] nl_BATCH_LOOP_acc_3_tmp;
  wire [7:0] STORE_LOOP_acc_2_tmp;
  wire [8:0] nl_STORE_LOOP_acc_2_tmp;
  wire [7:0] CALC_SOFTMAX_LOOP_acc_1_tmp;
  wire [8:0] nl_CALC_SOFTMAX_LOOP_acc_1_tmp;
  wire BATCH_LOOP_and_10_tmp;
  wire BATCH_LOOP_and_7_tmp;
  wire or_tmp_11;
  wire and_tmp_8;
  wire and_tmp_17;
  wire and_dcpl_29;
  wire and_dcpl_33;
  wire or_tmp_117;
  wire mux_tmp_151;
  wire and_dcpl_34;
  wire and_dcpl_36;
  wire and_dcpl_40;
  wire and_dcpl_43;
  wire and_dcpl_44;
  wire and_dcpl_45;
  wire mux_tmp_153;
  wire mux_tmp_154;
  wire or_dcpl_10;
  wire or_dcpl_30;
  wire or_dcpl_33;
  wire or_dcpl_39;
  wire mux_tmp_167;
  wire or_dcpl_40;
  wire or_dcpl_46;
  wire or_dcpl_47;
  wire or_dcpl_48;
  wire or_dcpl_49;
  wire and_dcpl_81;
  wire or_dcpl_50;
  wire and_dcpl_82;
  wire and_dcpl_84;
  wire mux_tmp_174;
  wire and_dcpl_92;
  wire and_dcpl_108;
  wire and_dcpl_110;
  wire nor_tmp_55;
  wire and_tmp_81;
  wire and_tmp_82;
  wire or_tmp_148;
  wire or_tmp_155;
  wire or_tmp_157;
  wire or_tmp_159;
  wire or_tmp_161;
  wire or_tmp_172;
  wire exit_BATCH_LOOP_lpi_1_dfm_mx1w0;
  wire CALC_SOFTMAX_LOOP_and_svs_1;
  wire CALC_SOFTMAX_LOOP_equal_tmp_2;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0;
  reg exitL_exit_CALC_SOFTMAX_LOOP_sva;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1;
  reg exit_BATCH_LOOP_lpi_1_dfm_st_3;
  reg BATCH_LOOP_stage_v_3;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0;
  reg exit_BATCH_LOOP_lpi_1_dfm_st_6;
  reg BATCH_LOOP_stage_v_6;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1;
  reg BATCH_LOOP_stage_v_7;
  wire CALC_SOFTMAX_LOOP_equal_tmp_3;
  wire CALC_SOFTMAX_LOOP_or_tmp_1;
  wire CALC_SOFTMAX_LOOP_and_10_ssc_1;
  wire CALC_SOFTMAX_LOOP_and_8_ssc_1;
  wire LOAD_LOOP_and_1_svs_1;
  wire [66:0] operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1;
  wire [73:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_sva_1_mx0w0;
  wire [74:0] nl_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_sva_1_mx0w0;
  reg BATCH_LOOP_stage_v_2;
  reg BATCH_LOOP_stage_0_3;
  reg BATCH_LOOP_stage_0_7;
  reg exit_BATCH_LOOP_lpi_1_dfm_st_7;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0;
  reg BATCH_LOOP_stage_v_5;
  reg BATCH_LOOP_stage_0_5;
  reg BATCH_LOOP_stage_0_6;
  reg BATCH_LOOP_stage_v_4;
  reg BATCH_LOOP_stage_0_4;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1;
  reg exit_BATCH_LOOP_lpi_1_dfm_st_2;
  reg exit_BATCH_LOOP_lpi_1_dfm_st_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0;
  reg BATCH_LOOP_stage_0;
  reg BATCH_LOOP_stage_v;
  reg CALC_SOFTMAX_LOOP_asn_itm;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1;
  reg CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_1;
  reg CALC_SOFTMAX_LOOP_asn_8_itm_1;
  reg CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_2;
  reg CALC_SOFTMAX_LOOP_asn_8_itm_2;
  reg BATCH_LOOP_stage_0_2;
  reg CALC_SOFTMAX_LOOP_asn_8_itm_3;
  reg CALC_SOFTMAX_LOOP_and_18_itm_3;
  reg CALC_SOFTMAX_LOOP_and_18_itm_2;
  reg LOAD_LOOP_and_1_svs_st_1;
  reg exit_BATCH_LOOP_sva_1_st_1;
  reg CALC_SOFTMAX_LOOP_asn_itm_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0;
  reg CALC_SOFTMAX_LOOP_asn_1_itm_1;
  wire [73:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_2;
  wire [73:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_mx1;
  wire and_210_m1c;
  wire asn_CALC_SOFTMAX_LOOP_i_7_0_lpi_1_6_0_nand_tmp;
  reg reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_cse;
  reg reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_cse;
  reg reg_dma_write_chnl_Push_mioi_iswt0_cse;
  reg reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_1_cse;
  wire CALC_SOFTMAX_LOOP_and_27_cse;
  wire and_413_cse;
  wire or_315_cse;
  wire or_323_cse;
  wire LOAD_LOOP_LOAD_LOOP_nor_1_cse;
  wire nand_93_cse;
  wire and_424_cse;
  wire nor_86_cse;
  wire mux_183_cse;
  wire mux_193_cse;
  wire mux_131_cse;
  wire mux_94_cse;
  wire mux_194_cse;
  reg [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d_reg;
  wire [66:0] operator_67_47_false_AC_TRN_AC_WRAP_mux_rmff;
  reg [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d_reg;
  wire [6:0] CALC_EXP_LOOP_i_mux_1_rmff;
  reg [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d_reg;
  wire [6:0] CALC_EXP_LOOP_i_mux_rmff;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff;
  wire and_241_rmff;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  wire and_245_rmff;
  wire and_243_rmff;
  wire [3:0] BATCH_LOOP_b_mux_rmff;
  wire BATCH_LOOP_BATCH_LOOP_or_11_rmff;
  wire LOAD_LOOP_LOAD_LOOP_or_rmff;
  wire [24:0] BATCH_LOOP_mux_rmff;
  wire BATCH_LOOP_BATCH_LOOP_or_12_rmff;
  wire [31:0] CALC_SOFTMAX_LOOP_mux_11_rmff;
  wire STORE_LOOP_STORE_LOOP_or_rmff;
  reg [93:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1;
  wire [93:0] operator_94_21_false_AC_TRN_AC_WRAP_rshift_itm;
  wire [72:0] operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm;
  reg [73:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1;
  reg [31:0] config_batch_sva;
  reg BATCH_LOOP_stage_v_1;
  reg exit_BATCH_LOOP_sva_1_st;
  reg LOAD_LOOP_and_1_svs_st;
  reg CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm;
  reg CALC_SOFTMAX_LOOP_and_18_itm;
  reg [93:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1_dfm_1;
  reg [73:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_sva_1_1;
  reg exit_BATCH_LOOP_sva_1_1;
  reg [73:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_1_1;
  reg [66:0] operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1_1;
  reg [6:0] CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_1;
  reg [6:0] CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_2;
  reg ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_itm_1;
  reg [6:0] CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_1;
  reg CALC_SOFTMAX_LOOP_and_18_itm_1;
  reg exit_BATCH_LOOP_lpi_1_dfm_st_4;
  reg exit_BATCH_LOOP_lpi_1_dfm_st_5;
  reg BATCH_LOOP_stage_0_1;
  reg [6:0] LOAD_LOOP_i_7_0_lpi_1_6_0;
  reg [6:0] CALC_EXP_LOOP_i_7_0_lpi_1_6_0;
  reg [6:0] SUM_EXP_LOOP_i_7_0_lpi_1_6_0;
  reg [6:0] CALC_SOFTMAX_LOOP_i_7_0_lpi_1_6_0;
  reg [3:0] BATCH_LOOP_b_4_0_sva_3_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1;
  reg lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_0;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_5_1_mx1w0;
  wire lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_5_0_mx1w0;
  wire CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_mx1w0;
  wire CALC_SOFTMAX_LOOP_and_18_itm_mx1w0;
  wire BATCH_LOOP_stage_0_mx1;
  wire CALC_SOFTMAX_LOOP_mux_10_mx1w0;
  wire BATCH_LOOP_BATCH_LOOP_or_10_cse_1;
  wire BATCH_LOOP_BATCH_LOOP_or_3_cse_1;
  wire BATCH_LOOP_BATCH_LOOP_or_2_cse_1;
  wire [18:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire [18:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire signed [19:0] nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1;
  wire CALC_SOFTMAX_LOOP_asn_65;
  wire [6:0] libraries_leading_sign_74_0_2abd7b3cff8691d03642c4ad577461acbee6_1;
  wire CALC_EXP_LOOP_i_and_2_rgt;
  wire dma_read_ctrl_write_reset_check_reset_nand_1_cse;
  wire CALC_SOFTMAX_LOOP_and_50_cse;
  wire CALC_SOFTMAX_LOOP_i_and_cse;
  wire CALC_SOFTMAX_LOOP_and_55_cse;
  wire CALC_SOFTMAX_LOOP_and_59_cse;
  wire CALC_SOFTMAX_LOOP_and_58_cse;
  wire BATCH_LOOP_and_18_cse;
  wire BATCH_LOOP_acc_1_itm_32_1;
  wire [18:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1;
  wire mux_209_cse;

  wire[0:0] or_242_nl;
  wire[0:0] or_248_nl;
  wire[0:0] or_249_nl;
  wire[24:0] BATCH_LOOP_acc_4_nl;
  wire[25:0] nl_BATCH_LOOP_acc_4_nl;
  wire[0:0] or_256_nl;
  wire[0:0] asn_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1_nand_nl;
  wire[0:0] and_152_nl;
  wire[0:0] and_153_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_i_and_3_nl;
  wire[0:0] and_167_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_or_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_and_48_nl;
  wire[0:0] mux_190_nl;
  wire[3:0] BATCH_LOOP_b_mux_2_nl;
  wire[0:0] BATCH_LOOP_b_and_nl;
  wire[0:0] BATCH_LOOP_mux1h_nl;
  wire[0:0] and_172_nl;
  wire[0:0] and_174_nl;
  wire[0:0] BATCH_LOOP_mux_47_nl;
  wire[0:0] asn_exitL_exit_CALC_SOFTMAX_LOOP_sva_nand_nl;
  wire[0:0] and_178_nl;
  wire[0:0] and_179_nl;
  wire[0:0] mux_196_nl;
  wire[0:0] and_426_nl;
  wire[0:0] mux_203_nl;
  wire[0:0] nor_63_nl;
  wire[0:0] mux_206_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] and_209_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_and_45_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_and_46_nl;
  wire[0:0] asn_LOAD_LOOP_i_7_0_lpi_1_6_0_nand_nl;
  wire[0:0] dma_read_ctrl_write_reset_check_ResetChecker_mux_nl;
  wire[0:0] BATCH_LOOP_mux_46_nl;
  wire[0:0] nor_94_nl;
  wire[0:0] BATCH_LOOP_mux_45_nl;
  wire[0:0] and_177_nl;
  wire[0:0] and_185_nl;
  wire[0:0] mux_192_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] and_186_nl;
  wire[0:0] BATCH_LOOP_mux_44_nl;
  wire[0:0] mux_195_nl;
  wire[0:0] nand_57_nl;
  wire[0:0] nand_58_nl;
  wire[0:0] BATCH_LOOP_mux_43_nl;
  wire[0:0] mux_200_nl;
  wire[0:0] nand_54_nl;
  wire[0:0] nand_55_nl;
  wire[0:0] BATCH_LOOP_mux_42_nl;
  wire[0:0] mux_201_nl;
  wire[0:0] BATCH_LOOP_mux_41_nl;
  wire[0:0] mux_202_nl;
  wire[0:0] and_214_nl;
  wire[0:0] and_55_nl;
  wire[0:0] CALC_SOFTMAX_LOOP_mux_34_nl;
  wire[0:0] and_160_nl;
  wire[0:0] and_163_nl;
  wire[0:0] or_187_nl;
  wire[32:0] BATCH_LOOP_acc_1_nl;
  wire[33:0] nl_BATCH_LOOP_acc_1_nl;
  wire[73:0] CALC_SOFTMAX_LOOP_mux_84_nl;
  wire[6:0] CALC_SOFTMAX_LOOP_mux_83_nl;
  wire[6:0] CALC_SOFTMAX_LOOP_mux_82_nl;
  wire[6:0] CALC_SOFTMAX_LOOP_mux_81_nl;
  wire[0:0] BATCH_LOOP_if_BATCH_LOOP_if_and_6_nl;
  wire[0:0] BATCH_LOOP_if_BATCH_LOOP_if_and_7_nl;
  wire[4:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_nl;
  wire[2:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_1_nl;
  wire[46:0] ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl;
  wire signed [47:0] nl_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl;
  wire[7:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_nl;
  wire[0:0] and_75_nl;
  wire[0:0] and_119_nl;
  wire[0:0] and_121_nl;
  wire[0:0] nand_61_nl;
  wire[0:0] mux_184_nl;
  wire[0:0] or_174_nl;
  wire[0:0] mux_189_nl;
  wire[0:0] mux_188_nl;
  wire[0:0] mux_187_nl;
  wire[0:0] mux_180_nl;
  wire[0:0] nor_69_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[10:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[9:0] ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl;
  wire [73:0] nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_a;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl
      = MUX_v_10_8_2(10'b1111111101, 10'b1100011001, 10'b1001100100, 10'b0111010000,
      10'b0101010100, 10'b0011101011, 10'b0010010001, 10'b0001000100, operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm[72:70]);
  assign nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_s2u_9_11(ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:10])
      + ({1'b1 , ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_1_nl});
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_a = {ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , (ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[9:0])
      , 53'b00000000000000000000000000000000000000000000000000000};
  wire [7:0] nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_s;
  assign nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_s = ({1'b1 , (~ libraries_leading_sign_74_0_2abd7b3cff8691d03642c4ad577461acbee6_1)})
      + 8'b00110111;
  wire[10:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[11:0] nl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl;
  wire[2:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_2_nl;
  wire[6:0] ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_3_nl;
  wire [20:0] nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_2_nl
      = MUX_v_3_4_2(3'b011, 3'b100, 3'b101, 3'b110, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1[11:10]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_3_nl
      = MUX_v_7_4_2(7'b1111110, 7'b1000000, 7'b0100110, 7'b0110111, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1[11:10]);
  assign nl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = conv_u2u_9_11(ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:10])
      + ({ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_2_nl
      , 1'b1 , ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_3_nl});
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl
      = nl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl[10:0];
  assign nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a = {ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_acc_nl
      , (ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[9:0])};
  wire [6:0] nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_s = ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1[18:12];
  wire [72:0] nl_operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg_a = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_sva_1_1[72:0];
  wire [31:0] nl_softmax_sysc_run_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat;
  assign nl_softmax_sysc_run_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat
      = {21'b000000000000000000000 , BATCH_LOOP_b_mux_rmff , 7'b0000000};
  wire [0:0] nl_softmax_sysc_run_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_oswt_unreg;
  assign nl_softmax_sysc_run_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_oswt_unreg
      = and_dcpl_29 & (fsm_output[2]);
  wire [0:0] nl_softmax_sysc_run_dma_read_chnl_Pop_mioi_inst_dma_read_chnl_Pop_mioi_oswt_unreg;
  assign nl_softmax_sysc_run_dma_read_chnl_Pop_mioi_inst_dma_read_chnl_Pop_mioi_oswt_unreg
      = and_dcpl_33 & (fsm_output[2]);
  wire [31:0] nl_softmax_sysc_run_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat;
  assign nl_softmax_sysc_run_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat
      = {BATCH_LOOP_mux_rmff , 7'b0000000};
  wire [0:0] nl_softmax_sysc_run_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_oswt_unreg;
  assign nl_softmax_sysc_run_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_oswt_unreg
      = and_dcpl_36 & (fsm_output[2]);
  wire [63:0] nl_softmax_sysc_run_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_m_rsc_dat;
  assign nl_softmax_sysc_run_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_m_rsc_dat
      = {32'b11011110101011011011111011101111 , CALC_SOFTMAX_LOOP_mux_11_rmff};
  wire [0:0] nl_softmax_sysc_run_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_oswt_unreg;
  assign nl_softmax_sysc_run_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_oswt_unreg
      = and_dcpl_44 & (fsm_output[2]);
  wire [0:0] nl_softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_inst_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg;
  assign nl_softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_inst_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg
      = mux_tmp_154 & BATCH_LOOP_stage_0_4 & ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1) & (~ exit_BATCH_LOOP_lpi_1_dfm_st_3)
      & BATCH_LOOP_stage_v_3 & (fsm_output[2]);
  wire [93:0] nl_softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp_inst_CALC_SOFTMAX_LOOP_mul_cmp_b_run;
  assign nl_softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp_inst_CALC_SOFTMAX_LOOP_mul_cmp_b_run
      = ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1;
  wire [0:0] nl_softmax_sysc_run_run_fsm_inst_CONFIG_LOOP_C_0_tr0;
  assign nl_softmax_sysc_run_run_fsm_inst_CONFIG_LOOP_C_0_tr0 = ~ conf_done;
  wire [0:0] nl_softmax_sysc_run_run_fsm_inst_BATCH_LOOP_C_0_tr0;
  assign nl_softmax_sysc_run_run_fsm_inst_BATCH_LOOP_C_0_tr0 = ~ BATCH_LOOP_nor_8_tmp;
  esp_acc_softmax_sysc_mgc_shift_br_v5 #(.width_a(32'sd74),
  .signd_a(32'sd0),
  .width_s(32'sd8),
  .width_z(32'sd94)) operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_a[73:0]),
      .s(nl_operator_94_21_false_AC_TRN_AC_WRAP_rshift_rg_s[7:0]),
      .z(operator_94_21_false_AC_TRN_AC_WRAP_rshift_itm)
    );
  esp_acc_softmax_sysc_mgc_shift_bl_v5 #(.width_a(32'sd21),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd67)) operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_a[20:0]),
      .s(nl_operator_67_47_false_AC_TRN_AC_WRAP_lshift_rg_s[6:0]),
      .z(operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1)
    );
  esp_acc_softmax_sysc_mgc_shift_l_v5 #(.width_a(32'sd73),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd73)) operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_operator_74_0_false_AC_TRN_AC_WRAP_lshift_rg_a[72:0]),
      .s(libraries_leading_sign_74_0_2abd7b3cff8691d03642c4ad577461acbee6_1),
      .z(operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm)
    );
  esp_acc_softmax_sysc_leading_sign_74_0  leading_sign_74_0_rg (
      .mantissa(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_sva_1_1),
      .rtn(libraries_leading_sign_74_0_2abd7b3cff8691d03642c4ad577461acbee6_1)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_dma_read_ctrl_Push_mioi softmax_sysc_run_dma_read_ctrl_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_ctrl_val(dma_read_ctrl_val),
      .dma_read_ctrl_rdy(dma_read_ctrl_rdy),
      .dma_read_ctrl_msg(dma_read_ctrl_msg),
      .run_wen(run_wen),
      .dma_read_ctrl_Push_mioi_m_index_rsc_dat(nl_softmax_sysc_run_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_m_index_rsc_dat[31:0]),
      .dma_read_ctrl_Push_mioi_oswt_unreg(nl_softmax_sysc_run_dma_read_ctrl_Push_mioi_inst_dma_read_ctrl_Push_mioi_oswt_unreg[0:0]),
      .dma_read_ctrl_Push_mioi_bawt(dma_read_ctrl_Push_mioi_bawt),
      .dma_read_ctrl_Push_mioi_iswt0(dma_read_ctrl_Push_mioi_iswt0),
      .run_wten(run_wten),
      .dma_read_ctrl_Push_mioi_wen_comp(dma_read_ctrl_Push_mioi_wen_comp),
      .dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct(BATCH_LOOP_BATCH_LOOP_or_11_rmff),
      .dma_read_ctrl_Push_mioi_iswt0_pff(or_tmp_155)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_dma_read_chnl_Pop_mioi softmax_sysc_run_dma_read_chnl_Pop_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_read_chnl_val(dma_read_chnl_val),
      .dma_read_chnl_rdy(dma_read_chnl_rdy),
      .dma_read_chnl_msg(dma_read_chnl_msg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .dma_read_chnl_Pop_mioi_oswt_unreg(nl_softmax_sysc_run_dma_read_chnl_Pop_mioi_inst_dma_read_chnl_Pop_mioi_oswt_unreg[0:0]),
      .dma_read_chnl_Pop_mioi_bawt(dma_read_chnl_Pop_mioi_bawt),
      .dma_read_chnl_Pop_mioi_iswt0(dma_read_chnl_Pop_mioi_iswt0),
      .dma_read_chnl_Pop_mioi_wen_comp(dma_read_chnl_Pop_mioi_wen_comp),
      .dma_read_chnl_Pop_mioi_return_rsc_z_mxwt(dma_read_chnl_Pop_mioi_return_rsc_z_mxwt),
      .dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_psct(LOAD_LOOP_LOAD_LOOP_or_rmff),
      .dma_read_chnl_Pop_mioi_iswt0_pff(or_tmp_157)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_dma_write_ctrl_Push_mioi softmax_sysc_run_dma_write_ctrl_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_ctrl_val(dma_write_ctrl_val),
      .dma_write_ctrl_rdy(dma_write_ctrl_rdy),
      .dma_write_ctrl_msg(dma_write_ctrl_msg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .dma_write_ctrl_Push_mioi_m_index_rsc_dat(nl_softmax_sysc_run_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_m_index_rsc_dat[31:0]),
      .dma_write_ctrl_Push_mioi_oswt_unreg(nl_softmax_sysc_run_dma_write_ctrl_Push_mioi_inst_dma_write_ctrl_Push_mioi_oswt_unreg[0:0]),
      .dma_write_ctrl_Push_mioi_bawt(dma_write_ctrl_Push_mioi_bawt),
      .dma_write_ctrl_Push_mioi_iswt0(dma_write_ctrl_Push_mioi_iswt0),
      .dma_write_ctrl_Push_mioi_wen_comp(dma_write_ctrl_Push_mioi_wen_comp),
      .dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct(BATCH_LOOP_BATCH_LOOP_or_12_rmff),
      .dma_write_ctrl_Push_mioi_iswt0_pff(or_tmp_159)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_dma_write_chnl_Push_mioi softmax_sysc_run_dma_write_chnl_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .dma_write_chnl_val(dma_write_chnl_val),
      .dma_write_chnl_rdy(dma_write_chnl_rdy),
      .dma_write_chnl_msg(dma_write_chnl_msg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .dma_write_chnl_Push_mioi_m_rsc_dat(nl_softmax_sysc_run_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_m_rsc_dat[63:0]),
      .dma_write_chnl_Push_mioi_oswt_unreg(nl_softmax_sysc_run_dma_write_chnl_Push_mioi_inst_dma_write_chnl_Push_mioi_oswt_unreg[0:0]),
      .dma_write_chnl_Push_mioi_bawt(dma_write_chnl_Push_mioi_bawt),
      .dma_write_chnl_Push_mioi_iswt0(reg_dma_write_chnl_Push_mioi_iswt0_cse),
      .dma_write_chnl_Push_mioi_wen_comp(dma_write_chnl_Push_mioi_wen_comp),
      .dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct(STORE_LOOP_STORE_LOOP_or_rmff),
      .dma_write_chnl_Push_mioi_iswt0_pff(or_tmp_161)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1
      softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg(nl_softmax_sysc_run_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_1_inst_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg[0:0]),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0(reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_cse),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_unreg_1(and_243_rmff),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1(reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_cse),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_pff(and_241_rmff),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_pff(and_245_rmff)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp_inst
      (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .CALC_SOFTMAX_LOOP_mul_cmp_oswt_unreg(or_tmp_161),
      .CALC_SOFTMAX_LOOP_mul_cmp_bawt(CALC_SOFTMAX_LOOP_mul_cmp_bawt),
      .CALC_SOFTMAX_LOOP_mul_cmp_iswt2(reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_1_cse),
      .CALC_SOFTMAX_LOOP_mul_cmp_a_run(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d_mxwt),
      .CALC_SOFTMAX_LOOP_mul_cmp_b_run(nl_softmax_sysc_run_CALC_SOFTMAX_LOOP_mul_cmp_inst_CALC_SOFTMAX_LOOP_mul_cmp_b_run[93:0]),
      .CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt(CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_staller softmax_sysc_run_staller_inst (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .dma_read_ctrl_Push_mioi_wen_comp(dma_read_ctrl_Push_mioi_wen_comp),
      .dma_read_chnl_Pop_mioi_wen_comp(dma_read_chnl_Pop_mioi_wen_comp),
      .dma_write_ctrl_Push_mioi_wen_comp(dma_write_ctrl_Push_mioi_wen_comp),
      .dma_write_chnl_Push_mioi_wen_comp(dma_write_chnl_Push_mioi_wen_comp)
    );
  esp_acc_softmax_sysc_softmax_sysc_run_run_fsm softmax_sysc_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .CONFIG_LOOP_C_0_tr0(nl_softmax_sysc_run_run_fsm_inst_CONFIG_LOOP_C_0_tr0[0:0]),
      .BATCH_LOOP_C_0_tr0(nl_softmax_sysc_run_run_fsm_inst_BATCH_LOOP_C_0_tr0[0:0])
    );
  assign and_241_rmff = mux_94_cse & and_413_cse & (~ exit_BATCH_LOOP_lpi_1_dfm_st_2)
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1) & (fsm_output[2]);
  assign and_243_rmff = mux_tmp_154 & BATCH_LOOP_stage_0_4 & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1
      & (~ exit_BATCH_LOOP_lpi_1_dfm_st_3) & BATCH_LOOP_stage_v_3 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0)
      & (fsm_output[2]);
  assign and_245_rmff = mux_94_cse & and_413_cse & (~ exit_BATCH_LOOP_lpi_1_dfm_st_2)
      & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0)
      & (fsm_output[2]);
  assign or_242_nl = (~ (fsm_output[2])) | (~((~(and_dcpl_43 & (~ dma_write_chnl_Push_mioi_bawt)
      & BATCH_LOOP_stage_v_7)) & CALC_SOFTMAX_LOOP_mul_cmp_bawt)) | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1)
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0 | exit_BATCH_LOOP_lpi_1_dfm_st_6
      | or_dcpl_10;
  assign CALC_SOFTMAX_LOOP_mux_11_rmff = MUX_v_32_2_2(CALC_SOFTMAX_LOOP_mul_cmp_z_mxwt,
      dma_write_chnl_Push_mioi_m_rsc_dat_31_0, or_242_nl);
  assign STORE_LOOP_STORE_LOOP_or_rmff = (dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct
      & (~(((~(CALC_SOFTMAX_LOOP_mul_cmp_bawt & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1))
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0 | exit_BATCH_LOOP_lpi_1_dfm_st_6
      | (~ BATCH_LOOP_stage_0_7) | (~ BATCH_LOOP_stage_v_6)) & and_dcpl_44 & (fsm_output[2]))))
      | or_tmp_161;
  assign CALC_EXP_LOOP_i_mux_rmff = MUX_v_7_2_2(CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_2,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d_reg,
      or_tmp_172);
  assign operator_67_47_false_AC_TRN_AC_WRAP_mux_rmff = MUX_v_67_2_2(operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d_reg,
      or_tmp_172);
  assign or_248_nl = (~ (fsm_output[2])) | (~ mux_94_cse) | nand_93_cse | exit_BATCH_LOOP_lpi_1_dfm_st_2
      | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1) | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0;
  assign CALC_EXP_LOOP_i_mux_1_rmff = MUX_v_7_2_2(CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_2,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d_reg,
      or_248_nl);
  assign or_249_nl = (~ (fsm_output[2])) | or_dcpl_30;
  assign BATCH_LOOP_b_mux_rmff = MUX_v_4_2_2(BATCH_LOOP_b_4_0_sva_3_0, dma_read_ctrl_Push_mioi_m_index_rsc_dat_10_7,
      or_249_nl);
  assign BATCH_LOOP_BATCH_LOOP_or_11_rmff = (dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct
      & (~(and_dcpl_29 & or_dcpl_30 & (fsm_output[2])))) | or_tmp_155;
  assign LOAD_LOOP_LOAD_LOOP_or_rmff = (dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_psct
      & (~(or_dcpl_33 & and_dcpl_33 & (fsm_output[2])))) | or_tmp_157;
  assign nl_BATCH_LOOP_acc_4_nl = (config_batch_sva[24:0]) + conv_u2u_4_25(BATCH_LOOP_b_4_0_sva_3_0);
  assign BATCH_LOOP_acc_4_nl = nl_BATCH_LOOP_acc_4_nl[24:0];
  assign or_256_nl = (~ (fsm_output[2])) | or_dcpl_39;
  assign BATCH_LOOP_mux_rmff = MUX_v_25_2_2(BATCH_LOOP_acc_4_nl, dma_write_ctrl_Push_mioi_m_index_rsc_dat_31_7,
      or_256_nl);
  assign BATCH_LOOP_BATCH_LOOP_or_12_rmff = (dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct
      & (~(or_dcpl_39 & and_dcpl_36 & (fsm_output[2])))) | or_tmp_159;
  assign CALC_SOFTMAX_LOOP_and_27_cse = run_wen & (fsm_output[2]);
  assign or_315_cse = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1 | exit_BATCH_LOOP_lpi_1_dfm_st_3;
  assign CALC_SOFTMAX_LOOP_and_50_cse = CALC_SOFTMAX_LOOP_and_27_cse & (~ exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign CALC_EXP_LOOP_i_and_2_rgt = exitL_exit_CALC_SOFTMAX_LOOP_sva & and_dcpl_34;
  assign CALC_SOFTMAX_LOOP_i_and_cse = CALC_SOFTMAX_LOOP_and_27_cse & BATCH_LOOP_and_10_tmp;
  assign CALC_SOFTMAX_LOOP_and_55_cse = CALC_SOFTMAX_LOOP_and_27_cse & mux_183_cse
      & BATCH_LOOP_and_10_tmp;
  assign mux_190_nl = MUX_s_1_2_2((~ BATCH_LOOP_stage_v), mux_tmp_174, BATCH_LOOP_and_10_tmp);
  assign dma_read_ctrl_write_reset_check_reset_nand_1_cse = ~(mux_190_nl & BATCH_LOOP_stage_0);
  assign CALC_SOFTMAX_LOOP_and_58_cse = run_wen & BATCH_LOOP_and_7_tmp;
  assign and_413_cse = BATCH_LOOP_stage_v_2 & BATCH_LOOP_stage_0_3;
  assign CALC_SOFTMAX_LOOP_and_59_cse = run_wen & ((~ BATCH_LOOP_stage_v_3) | exit_BATCH_LOOP_lpi_1_dfm_st_3
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1 | ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt)
      & and_tmp_8;
  assign nor_86_cse = ~(BATCH_LOOP_stage_v_6 | (~ or_tmp_11));
  assign mux_212_nl = MUX_s_1_2_2(LOAD_LOOP_and_1_svs_1, (~ CALC_SOFTMAX_LOOP_and_svs_1),
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1);
  assign mux_206_nl = MUX_s_1_2_2(mux_212_nl, LOAD_LOOP_and_1_svs_1, exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign and_210_m1c = mux_206_nl & BATCH_LOOP_and_10_tmp;
  assign mux_209_cse = MUX_s_1_2_2(nor_86_cse, or_tmp_11, or_323_cse);
  assign mux_214_nl = MUX_s_1_2_2(nor_86_cse, or_tmp_11, or_323_cse);
  assign mux_192_nl = MUX_s_1_2_2(nor_86_cse, mux_214_nl, BATCH_LOOP_stage_0_7);
  assign and_185_nl = BATCH_LOOP_stage_0_6 & mux_192_nl;
  assign mux_193_cse = MUX_s_1_2_2(mux_209_cse, and_185_nl, BATCH_LOOP_stage_v_5);
  assign and_186_nl = BATCH_LOOP_stage_0_5 & mux_193_cse;
  assign mux_194_cse = MUX_s_1_2_2(mux_209_cse, and_186_nl, BATCH_LOOP_stage_v_4);
  assign or_323_cse = CALC_SOFTMAX_LOOP_mul_cmp_bawt | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1)
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0 | exit_BATCH_LOOP_lpi_1_dfm_st_6;
  assign and_55_nl = or_315_cse & BATCH_LOOP_stage_0_4 & mux_194_cse;
  assign mux_94_cse = MUX_s_1_2_2(mux_209_cse, and_55_nl, BATCH_LOOP_stage_v_3);
  assign BATCH_LOOP_and_18_cse = run_wen & and_tmp_8;
  assign CALC_SOFTMAX_LOOP_mux_34_nl = MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0,
      (BATCH_LOOP_acc_3_tmp[4]), CALC_SOFTMAX_LOOP_and_10_ssc_1);
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_5_1_mx1w0 = CALC_SOFTMAX_LOOP_mux_34_nl
      | CALC_SOFTMAX_LOOP_and_8_ssc_1;
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_5_0_mx1w0 = (lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0
      & (~(CALC_SOFTMAX_LOOP_and_8_ssc_1 | CALC_SOFTMAX_LOOP_and_10_ssc_1))) | ((~
      LOAD_LOOP_and_1_svs_1) & CALC_SOFTMAX_LOOP_or_tmp_1);
  assign exit_BATCH_LOOP_lpi_1_dfm_mx1w0 = (~ BATCH_LOOP_acc_1_itm_32_1) & exitL_exit_CALC_SOFTMAX_LOOP_sva;
  assign and_160_nl = mux_94_cse & and_413_cse & (~ CALC_SOFTMAX_LOOP_asn_8_itm_2)
      & CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_2;
  assign and_163_nl = mux_94_cse & and_413_cse & (~(CALC_SOFTMAX_LOOP_asn_8_itm_2
      | CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_2));
  assign or_187_nl = (~ mux_94_cse) | nand_93_cse | CALC_SOFTMAX_LOOP_asn_8_itm_2;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_mx1
      = MUX1HOT_v_74_3_2(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_sva_1_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_1_1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1,
      {and_160_nl , and_163_nl , or_187_nl});
  assign nl_BATCH_LOOP_acc_1_nl = ({29'b10000000000000000000000000000 , BATCH_LOOP_b_4_0_sva_3_0})
      + conv_u2u_32_33(~ config_batch_sva) + 33'b000000000000000000000000000000001;
  assign BATCH_LOOP_acc_1_nl = nl_BATCH_LOOP_acc_1_nl[32:0];
  assign BATCH_LOOP_acc_1_itm_32_1 = readslicef_33_1_32(BATCH_LOOP_acc_1_nl);
  assign CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_mx1w0 = ~(CALC_SOFTMAX_LOOP_equal_tmp_2
      | CALC_SOFTMAX_LOOP_equal_tmp_3 | exit_BATCH_LOOP_lpi_1_dfm_mx1w0);
  assign CALC_SOFTMAX_LOOP_and_18_itm_mx1w0 = LOAD_LOOP_and_1_svs_1 & (~(CALC_SOFTMAX_LOOP_equal_tmp_2
      | CALC_SOFTMAX_LOOP_equal_tmp_3)) & (~ exit_BATCH_LOOP_lpi_1_dfm_mx1w0);
  assign BATCH_LOOP_stage_0_mx1 = BATCH_LOOP_stage_0 & (mux_tmp_174 | (~ BATCH_LOOP_and_10_tmp));
  assign CALC_SOFTMAX_LOOP_mux_10_mx1w0 = ~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_5_1_mx1w0
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_5_0_mx1w0);
  assign CALC_SOFTMAX_LOOP_mux_84_nl = MUX_v_74_2_2(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_mx1,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_2,
      CALC_SOFTMAX_LOOP_asn_1_itm_1);
  assign nl_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_sva_1_mx0w0
      = CALC_SOFTMAX_LOOP_mux_84_nl + conv_u2u_67_74(operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1);
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_sva_1_mx0w0
      = nl_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_sva_1_mx0w0[73:0];
  assign CALC_SOFTMAX_LOOP_equal_tmp_2 = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0);
  assign LOAD_LOOP_and_1_svs_1 = (LOAD_LOOP_acc_2_tmp[7]) & (CALC_EXP_LOOP_acc_1_tmp[7])
      & (SUM_EXP_LOOP_acc_2_tmp[7]);
  assign CALC_SOFTMAX_LOOP_mux_83_nl = MUX_v_7_2_2(LOAD_LOOP_i_7_0_lpi_1_6_0, (signext_7_1(~
      BATCH_LOOP_acc_1_itm_32_1)), exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign nl_LOAD_LOOP_acc_2_tmp = conv_u2u_7_8(CALC_SOFTMAX_LOOP_mux_83_nl) + 8'b00000001;
  assign LOAD_LOOP_acc_2_tmp = nl_LOAD_LOOP_acc_2_tmp[7:0];
  assign CALC_SOFTMAX_LOOP_mux_82_nl = MUX_v_7_2_2(CALC_EXP_LOOP_i_7_0_lpi_1_6_0,
      (signext_7_1(~ BATCH_LOOP_acc_1_itm_32_1)), exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign nl_CALC_EXP_LOOP_acc_1_tmp = conv_u2u_7_8(CALC_SOFTMAX_LOOP_mux_82_nl) +
      8'b00000001;
  assign CALC_EXP_LOOP_acc_1_tmp = nl_CALC_EXP_LOOP_acc_1_tmp[7:0];
  assign CALC_SOFTMAX_LOOP_mux_81_nl = MUX_v_7_2_2(SUM_EXP_LOOP_i_7_0_lpi_1_6_0,
      (signext_7_1(~ BATCH_LOOP_acc_1_itm_32_1)), exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign nl_SUM_EXP_LOOP_acc_2_tmp = conv_u2u_7_8(CALC_SOFTMAX_LOOP_mux_81_nl) +
      8'b00000001;
  assign SUM_EXP_LOOP_acc_2_tmp = nl_SUM_EXP_LOOP_acc_2_tmp[7:0];
  assign BATCH_LOOP_if_BATCH_LOOP_if_and_6_nl = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1
      & (~ BATCH_LOOP_acc_1_itm_32_1);
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0 = MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1,
      BATCH_LOOP_if_BATCH_LOOP_if_and_6_nl, exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign BATCH_LOOP_if_BATCH_LOOP_if_and_7_nl = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_0
      & (~ BATCH_LOOP_acc_1_itm_32_1);
  assign lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0 = MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_0,
      BATCH_LOOP_if_BATCH_LOOP_if_and_7_nl, exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign nl_BATCH_LOOP_acc_3_tmp = conv_u2u_4_5(BATCH_LOOP_b_4_0_sva_3_0) + 5'b00001;
  assign BATCH_LOOP_acc_3_tmp = nl_BATCH_LOOP_acc_3_tmp[4:0];
  assign CALC_SOFTMAX_LOOP_and_svs_1 = (CALC_SOFTMAX_LOOP_acc_1_tmp[7]) & (STORE_LOOP_acc_2_tmp[7]);
  assign nl_CALC_SOFTMAX_LOOP_acc_1_tmp = conv_u2u_7_8(CALC_SOFTMAX_LOOP_i_7_0_lpi_1_6_0)
      + 8'b00000001;
  assign CALC_SOFTMAX_LOOP_acc_1_tmp = nl_CALC_SOFTMAX_LOOP_acc_1_tmp[7:0];
  assign nl_STORE_LOOP_acc_2_tmp = conv_u2u_7_8(LOAD_LOOP_i_7_0_lpi_1_6_0) + 8'b00000001;
  assign STORE_LOOP_acc_2_tmp = nl_STORE_LOOP_acc_2_tmp[7:0];
  assign BATCH_LOOP_BATCH_LOOP_or_10_cse_1 = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_bawt
      | (~((~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1 | exit_BATCH_LOOP_lpi_1_dfm_st_3))
      & BATCH_LOOP_stage_v_3));
  assign BATCH_LOOP_BATCH_LOOP_or_3_cse_1 = CALC_SOFTMAX_LOOP_mul_cmp_bawt | (~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0) & (~ exit_BATCH_LOOP_lpi_1_dfm_st_6)
      & BATCH_LOOP_stage_v_6));
  assign BATCH_LOOP_BATCH_LOOP_or_2_cse_1 = dma_write_chnl_Push_mioi_bawt | (~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0) & (~ exit_BATCH_LOOP_lpi_1_dfm_st_7)
      & BATCH_LOOP_stage_v_7));
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_2
      = MUX_v_74_2_2(74'b00000000000000000000000000000000000000000000000000000000000000000000000000,
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_mx1,
      exit_BATCH_LOOP_sva_1_1);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_nl
      = MUX_v_5_4_2(5'b01100, 5'b01110, 5'b10001, 5'b10100, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1[11:10]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_1_nl
      = MUX_v_3_4_2(3'b010, 3'b110, 3'b001, 3'b101, ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1[11:10]);
  assign ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = conv_u2u_19_19(({ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_nl
      , 1'b0 , ac_math_ac_pow2_pwl_AC_TRN_33_7_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_output_pwl_mux_1_nl})
      * (ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1[9:0]));
  assign nl_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl
      = $signed((dma_read_chnl_Pop_mioi_return_rsc_z_mxwt)) * $signed(16'b0101110001010101);
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl
      = nl_ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl[46:0];
  assign ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_itm_46_28_1
      = readslicef_47_19_28(ac_math_ac_exp_pwl_0_AC_TRN_32_6_true_AC_TRN_AC_WRAP_67_47_AC_TRN_AC_WRAP_mul_nl);
  assign CALC_SOFTMAX_LOOP_equal_tmp_3 = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0
      & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0;
  assign CALC_SOFTMAX_LOOP_or_tmp_1 = (lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0)) | (~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0));
  assign CALC_SOFTMAX_LOOP_and_10_ssc_1 = CALC_SOFTMAX_LOOP_and_svs_1 & CALC_SOFTMAX_LOOP_equal_tmp_2;
  assign CALC_SOFTMAX_LOOP_and_8_ssc_1 = LOAD_LOOP_and_1_svs_1 & CALC_SOFTMAX_LOOP_or_tmp_1;
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_nl
      = MUX_v_8_8_2(8'b00011100, 8'b01001011, 8'b01101100, 8'b10000100, 8'b10010111,
      8'b10100110, 8'b10110011, 8'b10111100, operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm[72:70]);
  assign nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = $signed(({1'b1 , ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mux_nl}))
      * $signed(conv_u2s_10_11(operator_74_0_false_AC_TRN_AC_WRAP_lshift_itm[69:60]));
  assign ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1
      = nl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_pwl_mul_psp_sva_1[18:0];
  assign CALC_SOFTMAX_LOOP_asn_65 = CALC_SOFTMAX_LOOP_equal_tmp_2 & (~ exit_BATCH_LOOP_lpi_1_dfm_mx1w0);
  assign BATCH_LOOP_nor_8_tmp = ~((~(BATCH_LOOP_stage_v_7 & (dma_write_chnl_Push_mioi_bawt
      | (~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0)
      & (~ exit_BATCH_LOOP_lpi_1_dfm_st_7)))))) | BATCH_LOOP_stage_0_mx1 | BATCH_LOOP_stage_0_1
      | BATCH_LOOP_stage_0_2 | BATCH_LOOP_stage_0_3 | BATCH_LOOP_stage_0_4 | BATCH_LOOP_stage_0_5
      | BATCH_LOOP_stage_0_6 | BATCH_LOOP_stage_0_7);
  assign LOAD_LOOP_LOAD_LOOP_nor_1_cse = ~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1
      | exit_BATCH_LOOP_lpi_1_dfm_st_1);
  assign BATCH_LOOP_and_10_tmp = BATCH_LOOP_stage_v & (~(BATCH_LOOP_stage_v_1 & (~
      BATCH_LOOP_and_7_tmp))) & BATCH_LOOP_stage_0_1 & BATCH_LOOP_BATCH_LOOP_or_10_cse_1
      & BATCH_LOOP_BATCH_LOOP_or_3_cse_1 & BATCH_LOOP_BATCH_LOOP_or_2_cse_1;
  assign BATCH_LOOP_and_7_tmp = BATCH_LOOP_stage_v_1 & (~(BATCH_LOOP_stage_v_2 &
      or_dcpl_46)) & BATCH_LOOP_stage_0_2 & (dma_read_ctrl_Push_mioi_bawt | (~((~
      exit_BATCH_LOOP_sva_1_st_1) & CALC_SOFTMAX_LOOP_asn_itm_1))) & (dma_read_chnl_Pop_mioi_bawt
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1 | exit_BATCH_LOOP_lpi_1_dfm_st_1)
      & (dma_write_ctrl_Push_mioi_bawt | (~(LOAD_LOOP_and_1_svs_st_1 & ((lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1)) | (~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0))) & (~ exit_BATCH_LOOP_lpi_1_dfm_st_1))))
      & BATCH_LOOP_BATCH_LOOP_or_10_cse_1 & BATCH_LOOP_BATCH_LOOP_or_3_cse_1 & BATCH_LOOP_BATCH_LOOP_or_2_cse_1;
  assign or_tmp_11 = (~ BATCH_LOOP_stage_v_7) | dma_write_chnl_Push_mioi_bawt | exit_BATCH_LOOP_lpi_1_dfm_st_7
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0 | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1);
  assign and_tmp_8 = ((~ BATCH_LOOP_stage_v_6) | CALC_SOFTMAX_LOOP_mul_cmp_bawt |
      (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1) | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0
      | exit_BATCH_LOOP_lpi_1_dfm_st_6) & or_tmp_11;
  assign nand_93_cse = ~(BATCH_LOOP_stage_v_2 & BATCH_LOOP_stage_0_3);
  assign and_tmp_17 = or_323_cse & or_tmp_11;
  assign and_424_cse = BATCH_LOOP_stage_v_4 & BATCH_LOOP_stage_0_5;
  assign and_75_nl = BATCH_LOOP_stage_0_7 & and_tmp_17;
  assign mux_131_cse = MUX_s_1_2_2(or_tmp_11, and_75_nl, BATCH_LOOP_stage_v_6);
  assign and_dcpl_29 = CALC_SOFTMAX_LOOP_asn_itm_1 & (~ exit_BATCH_LOOP_sva_1_st_1)
      & BATCH_LOOP_and_7_tmp;
  assign and_dcpl_33 = LOAD_LOOP_LOAD_LOOP_nor_1_cse & BATCH_LOOP_and_7_tmp;
  assign or_tmp_117 = (~ CALC_SOFTMAX_LOOP_asn_itm) | BATCH_LOOP_acc_1_itm_32_1;
  assign mux_tmp_151 = MUX_s_1_2_2((~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1), or_tmp_117,
      exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign and_dcpl_34 = mux_tmp_151 & BATCH_LOOP_and_10_tmp;
  assign and_dcpl_36 = LOAD_LOOP_LOAD_LOOP_nor_1_cse & BATCH_LOOP_and_7_tmp & LOAD_LOOP_and_1_svs_st_1;
  assign and_dcpl_40 = mux_tmp_151 & (LOAD_LOOP_acc_2_tmp[7]) & (CALC_EXP_LOOP_acc_1_tmp[7])
      & (SUM_EXP_LOOP_acc_2_tmp[7]) & BATCH_LOOP_and_10_tmp;
  assign and_dcpl_43 = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1 & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0)
      & (~ exit_BATCH_LOOP_lpi_1_dfm_st_7);
  assign and_dcpl_44 = and_dcpl_43 & dma_write_chnl_Push_mioi_bawt & BATCH_LOOP_stage_v_7;
  assign and_dcpl_45 = BATCH_LOOP_stage_0_7 & BATCH_LOOP_stage_v_6;
  assign and_119_nl = BATCH_LOOP_stage_0_6 & mux_131_cse;
  assign mux_tmp_153 = MUX_s_1_2_2(and_tmp_8, and_119_nl, BATCH_LOOP_stage_v_5);
  assign and_121_nl = BATCH_LOOP_stage_0_5 & mux_tmp_153;
  assign mux_tmp_154 = MUX_s_1_2_2(and_tmp_8, and_121_nl, BATCH_LOOP_stage_v_4);
  assign or_dcpl_10 = ~(BATCH_LOOP_stage_0_7 & BATCH_LOOP_stage_v_6);
  assign or_dcpl_30 = ~(BATCH_LOOP_acc_1_itm_32_1 & CALC_SOFTMAX_LOOP_asn_itm & BATCH_LOOP_and_10_tmp);
  assign or_dcpl_33 = ~(mux_tmp_151 & BATCH_LOOP_and_10_tmp);
  assign or_dcpl_39 = ~(mux_tmp_151 & (LOAD_LOOP_acc_2_tmp[7]) & (CALC_EXP_LOOP_acc_1_tmp[7])
      & (SUM_EXP_LOOP_acc_2_tmp[7]) & BATCH_LOOP_and_10_tmp);
  assign mux_tmp_167 = or_tmp_117 & (SUM_EXP_LOOP_acc_2_tmp[7]) & (CALC_EXP_LOOP_acc_1_tmp[7])
      & (LOAD_LOOP_acc_2_tmp[7]);
  assign nand_61_nl = ~((BATCH_LOOP_acc_3_tmp[4]) & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1
      & (STORE_LOOP_acc_2_tmp[7]) & (CALC_SOFTMAX_LOOP_acc_1_tmp[7]));
  assign mux_183_cse = MUX_s_1_2_2(nand_61_nl, or_tmp_117, exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign or_174_nl = (~ exitL_exit_CALC_SOFTMAX_LOOP_sva) | (~ CALC_SOFTMAX_LOOP_asn_itm)
      | BATCH_LOOP_acc_1_itm_32_1;
  assign mux_184_nl = MUX_s_1_2_2(mux_183_cse, or_174_nl, lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_0);
  assign or_dcpl_40 = ~(mux_184_nl & BATCH_LOOP_and_10_tmp);
  assign or_dcpl_46 = (~ mux_94_cse) | nand_93_cse;
  assign or_dcpl_47 = ~(BATCH_LOOP_stage_0_6 & BATCH_LOOP_stage_v_5);
  assign or_dcpl_48 = (~ mux_131_cse) | or_dcpl_47;
  assign or_dcpl_49 = (~ and_tmp_17) | or_dcpl_10;
  assign and_dcpl_81 = (~ mux_tmp_151) & BATCH_LOOP_and_10_tmp;
  assign or_dcpl_50 = or_tmp_117 | (~ exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign and_dcpl_82 = or_dcpl_50 & BATCH_LOOP_and_10_tmp;
  assign and_dcpl_84 = (~ or_tmp_117) & exitL_exit_CALC_SOFTMAX_LOOP_sva & BATCH_LOOP_and_10_tmp;
  assign mux_tmp_174 = MUX_s_1_2_2(mux_183_cse, or_dcpl_50, lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_0);
  assign and_dcpl_92 = (~ mux_tmp_174) & BATCH_LOOP_and_10_tmp;
  assign and_dcpl_108 = BATCH_LOOP_stage_0_4 & BATCH_LOOP_stage_v_3;
  assign and_dcpl_110 = mux_tmp_154 & or_315_cse;
  assign nor_tmp_55 = BATCH_LOOP_stage_v_5 & BATCH_LOOP_stage_0_6;
  assign and_tmp_81 = nor_tmp_55 & mux_131_cse;
  assign and_tmp_82 = and_dcpl_45 & and_tmp_17;
  assign or_tmp_148 = dma_write_chnl_Push_mioi_bawt | exit_BATCH_LOOP_lpi_1_dfm_st_7
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0 | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1);
  assign or_tmp_155 = BATCH_LOOP_acc_1_itm_32_1 & CALC_SOFTMAX_LOOP_asn_itm & BATCH_LOOP_and_10_tmp
      & (fsm_output[2]);
  assign or_tmp_157 = and_dcpl_34 & (fsm_output[2]);
  assign or_tmp_159 = and_dcpl_40 & (fsm_output[2]);
  assign or_tmp_161 = or_tmp_11 & CALC_SOFTMAX_LOOP_mul_cmp_bawt & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1
      & (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0) & (~ exit_BATCH_LOOP_lpi_1_dfm_st_6)
      & and_dcpl_45 & (fsm_output[2]);
  assign or_tmp_172 = (~ (fsm_output[2])) | (~ mux_94_cse) | nand_93_cse | exit_BATCH_LOOP_lpi_1_dfm_st_2
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1;
  assign mux_187_nl = MUX_s_1_2_2(LOAD_LOOP_and_1_svs_1, (~ CALC_SOFTMAX_LOOP_and_svs_1),
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1);
  assign mux_188_nl = MUX_s_1_2_2(mux_187_nl, mux_tmp_167, exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign nor_69_nl = ~(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1 | (~ LOAD_LOOP_and_1_svs_1));
  assign mux_180_nl = MUX_s_1_2_2(nor_69_nl, mux_tmp_167, exitL_exit_CALC_SOFTMAX_LOOP_sva);
  assign mux_189_nl = MUX_s_1_2_2(mux_188_nl, mux_180_nl, lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_0);
  assign asn_CALC_SOFTMAX_LOOP_i_7_0_lpi_1_6_0_nand_tmp = ~(mux_189_nl & BATCH_LOOP_and_10_tmp);
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d
      = operator_67_47_false_AC_TRN_AC_WRAP_mux_rmff;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d
      = CALC_EXP_LOOP_i_mux_1_rmff;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d
      = CALC_EXP_LOOP_i_mux_rmff;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff;
  assign ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d
      = ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d_reg;
  always @(posedge clk) begin
    if ( ~ rst ) begin
      acc_done <= 1'b0;
    end
    else if ( run_wen & (((fsm_output[2]) & BATCH_LOOP_nor_8_tmp) | (fsm_output[5]))
        ) begin
      acc_done <= ~ (fsm_output[5]);
    end
  end
  always @(posedge clk) begin
    if ( run_wen ) begin
      dma_write_chnl_Push_mioi_m_rsc_dat_31_0 <= CALC_SOFTMAX_LOOP_mux_11_rmff;
      dma_write_chnl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct <= STORE_LOOP_STORE_LOOP_or_rmff;
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d_reg
          <= CALC_EXP_LOOP_i_mux_rmff;
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d_reg
          <= operator_67_47_false_AC_TRN_AC_WRAP_mux_rmff;
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d_reg
          <= CALC_EXP_LOOP_i_mux_1_rmff;
      dma_read_ctrl_Push_mioi_m_index_rsc_dat_10_7 <= BATCH_LOOP_b_mux_rmff;
      dma_read_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct <= BATCH_LOOP_BATCH_LOOP_or_11_rmff;
      dma_read_chnl_Pop_mioi_ccs_ccore_start_rsc_dat_run_psct <= LOAD_LOOP_LOAD_LOOP_or_rmff;
      dma_write_ctrl_Push_mioi_m_index_rsc_dat_31_7 <= BATCH_LOOP_mux_rmff;
      dma_write_ctrl_Push_mioi_ccs_ccore_start_rsc_dat_run_psct <= BATCH_LOOP_BATCH_LOOP_or_12_rmff;
      BATCH_LOOP_b_4_0_sva_3_0 <= MUX_v_4_2_2(4'b0000, BATCH_LOOP_b_mux_2_nl, (fsm_output[2]));
      config_batch_sva <= MUX_v_32_2_2(conf_info, config_batch_sva, fsm_output[2]);
      operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1_1 <= MUX_v_67_2_2(operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1_1,
          operator_67_47_false_AC_TRN_AC_WRAP_lshift_ncse_sva_1, BATCH_LOOP_and_7_tmp);
      CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_2 <= MUX1HOT_v_7_3_2(CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_1,
          CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_1, CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_2,
          {and_178_nl , and_179_nl , (~ BATCH_LOOP_and_7_tmp)});
      BATCH_LOOP_stage_v_1 <= ((BATCH_LOOP_stage_v_1 & (~ BATCH_LOOP_and_7_tmp))
          | BATCH_LOOP_and_10_tmp) & (fsm_output[2]);
      SUM_EXP_LOOP_i_7_0_lpi_1_6_0 <= MUX_v_7_2_2(SUM_EXP_LOOP_i_7_0_lpi_1_6_0, (SUM_EXP_LOOP_acc_2_tmp[6:0]),
          BATCH_LOOP_and_10_tmp);
      LOAD_LOOP_i_7_0_lpi_1_6_0 <= MUX1HOT_v_7_4_2((LOAD_LOOP_acc_2_tmp[6:0]), (signext_7_1(~
          LOAD_LOOP_and_1_svs_1)), (STORE_LOOP_acc_2_tmp[6:0]), LOAD_LOOP_i_7_0_lpi_1_6_0,
          {and_209_nl , CALC_SOFTMAX_LOOP_and_45_nl , CALC_SOFTMAX_LOOP_and_46_nl
          , asn_LOAD_LOOP_i_7_0_lpi_1_6_0_nand_nl});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      dma_read_ctrl_Push_mioi_iswt0 <= 1'b0;
      dma_read_chnl_Pop_mioi_iswt0 <= 1'b0;
      dma_write_ctrl_Push_mioi_iswt0 <= 1'b0;
      reg_dma_write_chnl_Push_mioi_iswt0_cse <= 1'b0;
      reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_cse
          <= 1'b0;
      reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_1_cse
          <= 1'b0;
      reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_cse
          <= 1'b0;
      BATCH_LOOP_stage_v <= 1'b0;
      BATCH_LOOP_stage_0 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm <= 1'b0;
      exitL_exit_CALC_SOFTMAX_LOOP_sva <= 1'b0;
      BATCH_LOOP_stage_v_2 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0 <= 1'b0;
      exit_BATCH_LOOP_lpi_1_dfm_st_2 <= 1'b0;
      BATCH_LOOP_stage_v_3 <= 1'b0;
      BATCH_LOOP_stage_v_4 <= 1'b0;
      BATCH_LOOP_stage_v_5 <= 1'b0;
      BATCH_LOOP_stage_v_6 <= 1'b0;
      BATCH_LOOP_stage_v_7 <= 1'b0;
      BATCH_LOOP_stage_0_1 <= 1'b0;
      BATCH_LOOP_stage_0_2 <= 1'b0;
      BATCH_LOOP_stage_0_3 <= 1'b0;
      BATCH_LOOP_stage_0_4 <= 1'b0;
      BATCH_LOOP_stage_0_5 <= 1'b0;
      BATCH_LOOP_stage_0_6 <= 1'b0;
      BATCH_LOOP_stage_0_7 <= 1'b0;
    end
    else if ( run_wen ) begin
      dma_read_ctrl_Push_mioi_iswt0 <= or_tmp_155;
      dma_read_chnl_Pop_mioi_iswt0 <= or_tmp_157;
      dma_write_ctrl_Push_mioi_iswt0 <= or_tmp_159;
      reg_dma_write_chnl_Push_mioi_iswt0_cse <= or_tmp_161;
      reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_cse
          <= and_241_rmff;
      reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_oswt_1_cse
          <= and_243_rmff;
      reg_ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_iswt0_1_cse
          <= and_245_rmff;
      BATCH_LOOP_stage_v <= ~((~(BATCH_LOOP_stage_v & (~((~(mux_tmp_174 & BATCH_LOOP_stage_0))
          & BATCH_LOOP_and_10_tmp)))) & dma_read_ctrl_write_reset_check_reset_nand_1_cse
          & (fsm_output[2]));
      BATCH_LOOP_stage_0 <= BATCH_LOOP_stage_0_mx1 | (~ (fsm_output[2]));
      CALC_SOFTMAX_LOOP_asn_itm <= BATCH_LOOP_mux1h_nl | (~ (fsm_output[2]));
      exitL_exit_CALC_SOFTMAX_LOOP_sva <= BATCH_LOOP_mux_47_nl | (~ (fsm_output[2]));
      BATCH_LOOP_stage_v_2 <= ((BATCH_LOOP_stage_v_2 & (~(mux_94_cse & and_413_cse)))
          | BATCH_LOOP_and_7_tmp) & (fsm_output[2]);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1, BATCH_LOOP_and_7_tmp);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0, BATCH_LOOP_and_7_tmp);
      exit_BATCH_LOOP_lpi_1_dfm_st_2 <= MUX_s_1_2_2(exit_BATCH_LOOP_lpi_1_dfm_st_2,
          exit_BATCH_LOOP_lpi_1_dfm_st_1, BATCH_LOOP_and_7_tmp);
      BATCH_LOOP_stage_v_3 <= ((BATCH_LOOP_stage_v_3 & (~(and_dcpl_110 & and_dcpl_108
          & nand_93_cse))) | (mux_94_cse & and_413_cse)) & (fsm_output[2]);
      BATCH_LOOP_stage_v_4 <= ((BATCH_LOOP_stage_v_4 & (~(mux_196_nl & and_424_cse)))
          | (and_dcpl_110 & and_dcpl_108)) & (fsm_output[2]);
      BATCH_LOOP_stage_v_5 <= ((BATCH_LOOP_stage_v_5 & (~(mux_131_cse & BATCH_LOOP_stage_0_6
          & (~(BATCH_LOOP_stage_0_5 & BATCH_LOOP_stage_v_4))))) | (mux_tmp_153 &
          and_424_cse)) & (fsm_output[2]);
      BATCH_LOOP_stage_v_6 <= ((BATCH_LOOP_stage_v_6 & (~(and_tmp_17 & and_dcpl_45
          & or_dcpl_47))) | and_tmp_81) & (fsm_output[2]);
      BATCH_LOOP_stage_v_7 <= ((BATCH_LOOP_stage_v_7 & (~ mux_203_nl)) | and_tmp_82)
          & (fsm_output[2]);
      BATCH_LOOP_stage_0_1 <= ~((~(dma_read_ctrl_write_reset_check_ResetChecker_mux_nl
          & (~ and_dcpl_92))) & (fsm_output[2]));
      BATCH_LOOP_stage_0_2 <= BATCH_LOOP_mux_46_nl & (fsm_output[2]);
      BATCH_LOOP_stage_0_3 <= BATCH_LOOP_mux_45_nl & (fsm_output[2]);
      BATCH_LOOP_stage_0_4 <= BATCH_LOOP_mux_44_nl & (fsm_output[2]);
      BATCH_LOOP_stage_0_5 <= BATCH_LOOP_mux_43_nl & (fsm_output[2]);
      BATCH_LOOP_stage_0_6 <= BATCH_LOOP_mux_42_nl & (fsm_output[2]);
      BATCH_LOOP_stage_0_7 <= BATCH_LOOP_mux_41_nl & (fsm_output[2]);
    end
  end
  always @(posedge clk) begin
    if ( CALC_SOFTMAX_LOOP_and_27_cse ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1
          <= MUX_v_94_2_2(ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1_dfm_1,
          ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1,
          asn_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1_nand_nl);
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1
          <= ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_mx1;
      CALC_EXP_LOOP_i_7_0_lpi_1_6_0 <= MUX1HOT_v_7_3_2((CALC_EXP_LOOP_acc_1_tmp[6:0]),
          CALC_EXP_LOOP_i_7_0_lpi_1_6_0, (signext_7_1(~ BATCH_LOOP_acc_1_itm_32_1)),
          {and_167_nl , CALC_SOFTMAX_LOOP_or_nl , CALC_SOFTMAX_LOOP_and_48_nl});
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1 <= 1'b0;
      exit_BATCH_LOOP_lpi_1_dfm_st_3 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0 <= 1'b0;
      exit_BATCH_LOOP_lpi_1_dfm_st_6 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0 <= 1'b0;
      exit_BATCH_LOOP_lpi_1_dfm_st_7 <= 1'b0;
      exit_BATCH_LOOP_sva_1_st_1 <= 1'b0;
      LOAD_LOOP_and_1_svs_st_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0 <= 1'b0;
      exit_BATCH_LOOP_lpi_1_dfm_st_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_itm_1 <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_27_cse ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_5_1_mx1w0,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1, or_dcpl_40);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_1,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1, or_dcpl_46);
      exit_BATCH_LOOP_lpi_1_dfm_st_3 <= MUX_s_1_2_2(exit_BATCH_LOOP_lpi_1_dfm_st_2,
          exit_BATCH_LOOP_lpi_1_dfm_st_3, or_dcpl_46);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1, or_dcpl_48);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_0,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0, or_dcpl_48);
      exit_BATCH_LOOP_lpi_1_dfm_st_6 <= MUX_s_1_2_2(exit_BATCH_LOOP_lpi_1_dfm_st_5,
          exit_BATCH_LOOP_lpi_1_dfm_st_6, or_dcpl_48);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_1,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_1, or_dcpl_49);
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0 <= MUX_s_1_2_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_6_0,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_7_0, or_dcpl_49);
      exit_BATCH_LOOP_lpi_1_dfm_st_7 <= MUX_s_1_2_2(exit_BATCH_LOOP_lpi_1_dfm_st_6,
          exit_BATCH_LOOP_lpi_1_dfm_st_7, or_dcpl_49);
      exit_BATCH_LOOP_sva_1_st_1 <= MUX1HOT_s_1_3_2((~ BATCH_LOOP_acc_1_itm_32_1),
          exit_BATCH_LOOP_sva_1_st, exit_BATCH_LOOP_sva_1_st_1, {and_152_nl , and_153_nl
          , (~ BATCH_LOOP_and_10_tmp)});
      LOAD_LOOP_and_1_svs_st_1 <= MUX1HOT_s_1_3_2(LOAD_LOOP_and_1_svs_1, LOAD_LOOP_and_1_svs_st,
          LOAD_LOOP_and_1_svs_st_1, {and_dcpl_34 , and_dcpl_81 , (~ BATCH_LOOP_and_10_tmp)});
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1 <= MUX1HOT_s_1_3_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_1_mx0,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1, lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1,
          {and_dcpl_82 , and_dcpl_84 , (~ BATCH_LOOP_and_10_tmp)});
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0 <= MUX1HOT_s_1_3_2(lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_0_mx0,
          lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_0, lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_0,
          {and_dcpl_82 , and_dcpl_84 , (~ BATCH_LOOP_and_10_tmp)});
      exit_BATCH_LOOP_lpi_1_dfm_st_1 <= MUX_s_1_2_2(exit_BATCH_LOOP_lpi_1_dfm_st_1,
          exit_BATCH_LOOP_lpi_1_dfm_mx1w0, BATCH_LOOP_and_10_tmp);
      CALC_SOFTMAX_LOOP_asn_itm_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_asn_itm_1, CALC_SOFTMAX_LOOP_asn_itm,
          BATCH_LOOP_and_10_tmp);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_0 <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_27_cse & (~ or_dcpl_40) ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_5_0_mx1w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      LOAD_LOOP_and_1_svs_st <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_27_cse & (~ or_dcpl_33) ) begin
      LOAD_LOOP_and_1_svs_st <= LOAD_LOOP_and_1_svs_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_0 <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_50_cse ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_0;
    end
  end
  always @(posedge clk) begin
    if ( CALC_SOFTMAX_LOOP_and_27_cse & (((~ exitL_exit_CALC_SOFTMAX_LOOP_sva) &
        and_dcpl_34) | and_dcpl_81 | CALC_EXP_LOOP_i_and_2_rgt) ) begin
      CALC_EXP_LOOP_i_slc_CALC_EXP_LOOP_i_7_0_6_0_1_itm_1 <= MUX_v_7_2_2(CALC_EXP_LOOP_i_7_0_lpi_1_6_0,
          (signext_7_1(~ BATCH_LOOP_acc_1_itm_32_1)), CALC_EXP_LOOP_i_and_2_rgt);
    end
  end
  always @(posedge clk) begin
    if ( CALC_SOFTMAX_LOOP_i_and_cse ) begin
      CALC_SOFTMAX_LOOP_i_slc_CALC_SOFTMAX_LOOP_i_7_0_6_0_itm_1 <= CALC_SOFTMAX_LOOP_i_7_0_lpi_1_6_0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_asn_8_itm_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_1_itm_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_1 <= 1'b0;
      CALC_SOFTMAX_LOOP_and_18_itm_1 <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_i_and_cse ) begin
      CALC_SOFTMAX_LOOP_asn_8_itm_1 <= ((BATCH_LOOP_acc_3_tmp[4]) & CALC_SOFTMAX_LOOP_and_svs_1
          & CALC_SOFTMAX_LOOP_equal_tmp_2) | exit_BATCH_LOOP_lpi_1_dfm_mx1w0;
      CALC_SOFTMAX_LOOP_asn_1_itm_1 <= exitL_exit_CALC_SOFTMAX_LOOP_sva;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_mx1w0,
          CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm, and_dcpl_92);
      CALC_SOFTMAX_LOOP_and_18_itm_1 <= MUX_s_1_2_2(CALC_SOFTMAX_LOOP_and_18_itm_mx1w0,
          CALC_SOFTMAX_LOOP_and_18_itm, and_dcpl_92);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_BATCH_LOOP_sva_1_1 <= 1'b0;
    end
    else if ( run_wen & BATCH_LOOP_and_10_tmp & (fsm_output[2]) ) begin
      exit_BATCH_LOOP_sva_1_1 <= ~ BATCH_LOOP_acc_1_itm_32_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm <= 1'b0;
      CALC_SOFTMAX_LOOP_and_18_itm <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_55_cse ) begin
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm <= CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_mx1w0;
      CALC_SOFTMAX_LOOP_and_18_itm <= CALC_SOFTMAX_LOOP_and_18_itm_mx1w0;
    end
  end
  always @(posedge clk) begin
    if ( CALC_SOFTMAX_LOOP_and_27_cse & (~ asn_CALC_SOFTMAX_LOOP_i_7_0_lpi_1_6_0_nand_tmp)
        ) begin
      CALC_SOFTMAX_LOOP_i_7_0_lpi_1_6_0 <= MUX_v_7_2_2((signext_7_1(~ LOAD_LOOP_and_1_svs_1)),
          (CALC_SOFTMAX_LOOP_acc_1_tmp[6:0]), CALC_SOFTMAX_LOOP_i_and_3_nl);
    end
  end
  always @(posedge clk) begin
    if ( CALC_SOFTMAX_LOOP_and_58_cse ) begin
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_1_1
          <= MUX_v_74_2_2(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_dfm_2,
          ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_lpi_1_mx1,
          and_214_nl);
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_sva_1_1
          <= ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_sva_1_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      CALC_SOFTMAX_LOOP_asn_8_itm_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_2 <= 1'b0;
      CALC_SOFTMAX_LOOP_and_18_itm_2 <= 1'b0;
      ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_itm_1
          <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_58_cse ) begin
      CALC_SOFTMAX_LOOP_asn_8_itm_2 <= CALC_SOFTMAX_LOOP_asn_8_itm_1;
      CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_2 <= CALC_SOFTMAX_LOOP_CALC_SOFTMAX_LOOP_nor_2_itm_1;
      CALC_SOFTMAX_LOOP_and_18_itm_2 <= CALC_SOFTMAX_LOOP_and_18_itm_1;
      ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_itm_1
          <= ~((ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_sum_exp_sva_1_mx0w0!=74'b00000000000000000000000000000000000000000000000000000000000000000000000000));
    end
  end
  always @(posedge clk) begin
    if ( CALC_SOFTMAX_LOOP_and_59_cse ) begin
      ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1_dfm_1
          <= MUX_v_94_2_2(operator_94_21_false_AC_TRN_AC_WRAP_rshift_itm, 94'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
          ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_ac_math_ac_normalize_74_54_false_AC_TRN_AC_WRAP_expret_nor_itm_1);
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0 <= 1'b0;
      CALC_SOFTMAX_LOOP_asn_8_itm_3 <= 1'b0;
      CALC_SOFTMAX_LOOP_and_18_itm_3 <= 1'b0;
    end
    else if ( CALC_SOFTMAX_LOOP_and_59_cse ) begin
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_2_0;
      CALC_SOFTMAX_LOOP_asn_8_itm_3 <= CALC_SOFTMAX_LOOP_asn_8_itm_2;
      CALC_SOFTMAX_LOOP_and_18_itm_3 <= CALC_SOFTMAX_LOOP_and_18_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_BATCH_LOOP_sva_1_st <= 1'b0;
    end
    else if ( run_wen & CALC_SOFTMAX_LOOP_asn_itm & BATCH_LOOP_and_10_tmp ) begin
      exit_BATCH_LOOP_sva_1_st <= ~ BATCH_LOOP_acc_1_itm_32_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ rst ) begin
      exit_BATCH_LOOP_lpi_1_dfm_st_5 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_0 <= 1'b0;
      exit_BATCH_LOOP_lpi_1_dfm_st_4 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1 <= 1'b0;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0 <= 1'b0;
    end
    else if ( BATCH_LOOP_and_18_cse ) begin
      exit_BATCH_LOOP_lpi_1_dfm_st_5 <= exit_BATCH_LOOP_lpi_1_dfm_st_4;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_5_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0;
      exit_BATCH_LOOP_lpi_1_dfm_st_4 <= exit_BATCH_LOOP_lpi_1_dfm_st_3;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_1 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_1;
      lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_4_0 <= lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_3_0;
    end
  end
  assign BATCH_LOOP_b_and_nl = ((~((CALC_SOFTMAX_LOOP_acc_1_tmp[7]) & (STORE_LOOP_acc_2_tmp[7])))
      | (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1) | (BATCH_LOOP_acc_3_tmp[4]) | exitL_exit_CALC_SOFTMAX_LOOP_sva
      | lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_0 | (~ BATCH_LOOP_and_10_tmp)) & (fsm_output[2]);
  assign BATCH_LOOP_b_mux_2_nl = MUX_v_4_2_2((BATCH_LOOP_acc_3_tmp[3:0]), BATCH_LOOP_b_4_0_sva_3_0,
      BATCH_LOOP_b_and_nl);
  assign and_172_nl = mux_tmp_174 & BATCH_LOOP_stage_0 & BATCH_LOOP_and_10_tmp;
  assign and_174_nl = (~ BATCH_LOOP_stage_v) & BATCH_LOOP_stage_0;
  assign BATCH_LOOP_mux1h_nl = MUX1HOT_s_1_3_2(CALC_SOFTMAX_LOOP_mux_10_mx1w0, exitL_exit_CALC_SOFTMAX_LOOP_sva,
      CALC_SOFTMAX_LOOP_asn_itm, {and_172_nl , and_174_nl , dma_read_ctrl_write_reset_check_reset_nand_1_cse});
  assign asn_exitL_exit_CALC_SOFTMAX_LOOP_sva_nand_nl = ~(mux_tmp_174 & BATCH_LOOP_and_10_tmp);
  assign BATCH_LOOP_mux_47_nl = MUX_s_1_2_2(CALC_SOFTMAX_LOOP_mux_10_mx1w0, exitL_exit_CALC_SOFTMAX_LOOP_sva,
      asn_exitL_exit_CALC_SOFTMAX_LOOP_sva_nand_nl);
  assign and_178_nl = (~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1) & BATCH_LOOP_and_7_tmp;
  assign and_179_nl = lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_dfm_1_st_1_1 & BATCH_LOOP_and_7_tmp;
  assign and_426_nl = (~(or_315_cse & BATCH_LOOP_stage_0_4)) & mux_tmp_153;
  assign mux_196_nl = MUX_s_1_2_2(mux_tmp_153, and_426_nl, BATCH_LOOP_stage_v_3);
  assign nor_63_nl = ~(or_323_cse | (~ or_tmp_148));
  assign mux_203_nl = MUX_s_1_2_2(or_tmp_148, nor_63_nl, and_dcpl_45);
  assign and_209_nl = (~(LOAD_LOOP_and_1_svs_1 | (~((~ lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1)
      | exitL_exit_CALC_SOFTMAX_LOOP_sva)))) & BATCH_LOOP_and_10_tmp;
  assign CALC_SOFTMAX_LOOP_and_45_nl = (~ CALC_SOFTMAX_LOOP_asn_65) & and_210_m1c;
  assign CALC_SOFTMAX_LOOP_and_46_nl = CALC_SOFTMAX_LOOP_asn_65 & and_210_m1c;
  assign asn_LOAD_LOOP_i_7_0_lpi_1_6_0_nand_nl = ~((~(CALC_SOFTMAX_LOOP_and_svs_1
      & lfst_exit_CALC_SOFTMAX_LOOP_lpi_1_1 & (~ exitL_exit_CALC_SOFTMAX_LOOP_sva)))
      & BATCH_LOOP_and_10_tmp);
  assign dma_read_ctrl_write_reset_check_ResetChecker_mux_nl = MUX_s_1_2_2(BATCH_LOOP_stage_0_1,
      BATCH_LOOP_stage_0, BATCH_LOOP_and_10_tmp);
  assign nor_94_nl = ~(BATCH_LOOP_and_7_tmp | BATCH_LOOP_and_10_tmp);
  assign BATCH_LOOP_mux_46_nl = MUX_s_1_2_2(BATCH_LOOP_stage_0_1, BATCH_LOOP_stage_0_2,
      nor_94_nl);
  assign and_177_nl = or_dcpl_46 & (~ BATCH_LOOP_and_7_tmp);
  assign BATCH_LOOP_mux_45_nl = MUX_s_1_2_2(BATCH_LOOP_stage_0_2, BATCH_LOOP_stage_0_3,
      and_177_nl);
  assign nand_57_nl = ~(BATCH_LOOP_stage_v_2 & BATCH_LOOP_stage_0_3 & mux_209_cse);
  assign nand_58_nl = ~(or_315_cse & BATCH_LOOP_stage_0_4 & mux_194_cse);
  assign mux_195_nl = MUX_s_1_2_2(nand_57_nl, nand_58_nl, BATCH_LOOP_stage_v_3);
  assign BATCH_LOOP_mux_44_nl = MUX_s_1_2_2(BATCH_LOOP_stage_0_3, BATCH_LOOP_stage_0_4,
      mux_195_nl);
  assign nand_54_nl = ~(or_315_cse & BATCH_LOOP_stage_v_3 & BATCH_LOOP_stage_0_4
      & mux_209_cse);
  assign nand_55_nl = ~(BATCH_LOOP_stage_0_5 & mux_193_cse);
  assign mux_200_nl = MUX_s_1_2_2(nand_54_nl, nand_55_nl, BATCH_LOOP_stage_v_4);
  assign BATCH_LOOP_mux_43_nl = MUX_s_1_2_2(BATCH_LOOP_stage_0_4, BATCH_LOOP_stage_0_5,
      mux_200_nl);
  assign mux_201_nl = MUX_s_1_2_2(and_tmp_81, mux_tmp_153, and_424_cse);
  assign BATCH_LOOP_mux_42_nl = MUX_s_1_2_2(BATCH_LOOP_stage_0_6, BATCH_LOOP_stage_0_5,
      mux_201_nl);
  assign mux_202_nl = MUX_s_1_2_2(and_tmp_82, mux_131_cse, nor_tmp_55);
  assign BATCH_LOOP_mux_41_nl = MUX_s_1_2_2(BATCH_LOOP_stage_0_7, BATCH_LOOP_stage_0_6,
      mux_202_nl);
  assign asn_ac_math_ac_reciprocal_pwl_AC_TRN_74_54_false_AC_TRN_AC_WRAP_94_21_false_AC_TRN_AC_WRAP_output_temp_lpi_1_nand_nl
      = ~(mux_tmp_154 & or_315_cse & BATCH_LOOP_stage_0_4 & BATCH_LOOP_stage_v_3
      & (~ CALC_SOFTMAX_LOOP_asn_8_itm_3) & CALC_SOFTMAX_LOOP_and_18_itm_3);
  assign and_152_nl = CALC_SOFTMAX_LOOP_asn_itm & BATCH_LOOP_and_10_tmp;
  assign and_153_nl = (~ CALC_SOFTMAX_LOOP_asn_itm) & BATCH_LOOP_and_10_tmp;
  assign and_167_nl = mux_tmp_151 & (~ LOAD_LOOP_and_1_svs_1) & BATCH_LOOP_and_10_tmp;
  assign CALC_SOFTMAX_LOOP_or_nl = ((~ exitL_exit_CALC_SOFTMAX_LOOP_sva) & and_dcpl_40)
      | or_dcpl_33;
  assign CALC_SOFTMAX_LOOP_and_48_nl = exitL_exit_CALC_SOFTMAX_LOOP_sva & and_dcpl_40;
  assign CALC_SOFTMAX_LOOP_i_and_3_nl = CALC_SOFTMAX_LOOP_asn_65 & (~ asn_CALC_SOFTMAX_LOOP_i_7_0_lpi_1_6_0_nand_tmp);
  assign and_214_nl = BATCH_LOOP_and_7_tmp & (~ CALC_SOFTMAX_LOOP_asn_1_itm_1);

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [73:0] MUX1HOT_v_74_3_2;
    input [73:0] input_2;
    input [73:0] input_1;
    input [73:0] input_0;
    input [2:0] sel;
    reg [73:0] result;
  begin
    result = input_0 & {74{sel[0]}};
    result = result | ( input_1 & {74{sel[1]}});
    result = result | ( input_2 & {74{sel[2]}});
    MUX1HOT_v_74_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_4_2;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [3:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    result = result | ( input_3 & {7{sel[3]}});
    MUX1HOT_v_7_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_8_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [9:0] input_2;
    input [9:0] input_3;
    input [9:0] input_4;
    input [9:0] input_5;
    input [9:0] input_6;
    input [9:0] input_7;
    input [2:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_10_8_2 = result;
  end
  endfunction


  function automatic [24:0] MUX_v_25_2_2;
    input [24:0] input_0;
    input [24:0] input_1;
    input [0:0] sel;
    reg [24:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_25_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_4_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [1:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_3_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_4_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [4:0] input_2;
    input [4:0] input_3;
    input [1:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_5_4_2 = result;
  end
  endfunction


  function automatic [66:0] MUX_v_67_2_2;
    input [66:0] input_0;
    input [66:0] input_1;
    input [0:0] sel;
    reg [66:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_67_2_2 = result;
  end
  endfunction


  function automatic [73:0] MUX_v_74_2_2;
    input [73:0] input_0;
    input [73:0] input_1;
    input [0:0] sel;
    reg [73:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_74_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_4_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [6:0] input_2;
    input [6:0] input_3;
    input [1:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_7_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_8_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2 = result;
  end
  endfunction


  function automatic [93:0] MUX_v_94_2_2;
    input [93:0] input_0;
    input [93:0] input_1;
    input [0:0] sel;
    reg [93:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_94_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [18:0] readslicef_47_19_28;
    input [46:0] vector;
    reg [46:0] tmp;
  begin
    tmp = vector >> 28;
    readslicef_47_19_28 = tmp[18:0];
  end
  endfunction


  function automatic [6:0] signext_7_1;
    input [0:0] vector;
  begin
    signext_7_1= {{6{vector[0]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_s2u_9_11 = {{2{vector[8]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function automatic [24:0] conv_u2u_4_25 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_25 = {{21{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_9_11 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_11 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [18:0] conv_u2u_19_19 ;
    input [18:0]  vector ;
  begin
    conv_u2u_19_19 = vector;
  end
  endfunction


  function automatic [32:0] conv_u2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_33 = {1'b0, vector};
  end
  endfunction


  function automatic [73:0] conv_u2u_67_74 ;
    input [66:0]  vector ;
  begin
    conv_u2u_67_74 = {{7{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    softmax_sysc_basic_fx32_dma64
// ------------------------------------------------------------------


module softmax_sysc_basic_fx32_dma64 (
  clk, rst, conf_info, conf_done, acc_done, debug, dma_read_ctrl_val, dma_read_ctrl_rdy,
      dma_read_ctrl_msg, dma_write_ctrl_val, dma_write_ctrl_rdy, dma_write_ctrl_msg,
      dma_read_chnl_val, dma_read_chnl_rdy, dma_read_chnl_msg, dma_write_chnl_val,
      dma_write_chnl_rdy, dma_write_chnl_msg
);
  input clk;
  input rst;
  input [31:0] conf_info;
  input conf_done;
  output acc_done;
  output [31:0] debug;
  output dma_read_ctrl_val;
  input dma_read_ctrl_rdy;
  output [66:0] dma_read_ctrl_msg;
  output dma_write_ctrl_val;
  input dma_write_ctrl_rdy;
  output [66:0] dma_write_ctrl_msg;
  input dma_read_chnl_val;
  output dma_read_chnl_rdy;
  input [63:0] dma_read_chnl_msg;
  output dma_write_chnl_val;
  input dma_write_chnl_rdy;
  output [63:0] dma_write_chnl_msg;


  // Interconnect Declarations
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_clken;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_q;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_radr;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_we;
  wire [66:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_d;
  wire [6:0] ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wadr;
  wire ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  BLOCK_1R1W_RBW #(.addr_width(32'sd7),
  .data_width(32'sd67),
  .depth(32'sd128),
  .latency(32'sd1)) ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_comp
      (
      .clk(clk),
      .clken(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_clken),
      .d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_d),
      .q(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_q),
      .radr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_radr),
      .wadr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wadr),
      .we(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_we)
    );
  esp_acc_softmax_sysc_softmax_sysc_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_en_12_7_67_128_128_67_1_gen
      ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci
      (
      .clken(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_clken),
      .q(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_q),
      .radr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_radr),
      .we(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_we),
      .d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_d),
      .wadr(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsc_wadr),
      .clken_d(1'b1),
      .d_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d),
      .q_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d),
      .radr_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d),
      .wadr_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d),
      .we_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d)
    );
  esp_acc_softmax_sysc_softmax_sysc_run softmax_sysc_run_inst (
      .clk(clk),
      .rst(rst),
      .conf_info(conf_info),
      .conf_done(conf_done),
      .acc_done(acc_done),
      .dma_read_ctrl_val(dma_read_ctrl_val),
      .dma_read_ctrl_rdy(dma_read_ctrl_rdy),
      .dma_read_ctrl_msg(dma_read_ctrl_msg),
      .dma_write_ctrl_val(dma_write_ctrl_val),
      .dma_write_ctrl_rdy(dma_write_ctrl_rdy),
      .dma_write_ctrl_msg(dma_write_ctrl_msg),
      .dma_read_chnl_val(dma_read_chnl_val),
      .dma_read_chnl_rdy(dma_read_chnl_rdy),
      .dma_read_chnl_msg(dma_read_chnl_msg),
      .dma_write_chnl_val(dma_write_chnl_val),
      .dma_write_chnl_rdy(dma_write_chnl_rdy),
      .dma_write_chnl_msg(dma_write_chnl_msg),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_d_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_q_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_radr_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_wadr_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_readA_r_ram_ir_internal_RMASK_B_d),
      .ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_pff(ac_math_ac_softmax_pwl_AC_TRN_false_0_0_AC_TRN_AC_WRAP_false_0_0_AC_TRN_AC_WRAP_128U_32_6_true_AC_TRN_AC_WRAP_32_2_AC_TRN_AC_WRAP_exp_arr_rsci_we_d_iff)
    );
  assign debug = 32'b00000000000000000000000000000000;
endmodule



